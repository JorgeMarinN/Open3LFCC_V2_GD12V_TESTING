magic
tech sky130A
timestamp 1675430904
<< error_p >>
rect 507 607 610 663
rect 497 575 1075 607
rect 81 553 1075 575
rect 345 550 385 553
rect 497 550 1075 553
rect -25 205 -3 469
rect 156 447 160 550
rect 787 547 1063 550
rect -25 160 0 205
rect -25 156 156 160
rect -25 117 160 156
rect -25 43 -3 117
rect 0 43 160 117
rect -113 0 160 43
rect -113 -113 43 0
rect 147 -21 205 0
<< pwell >>
rect 0 0 1175 550
<< mvnmos >>
rect 81 500 519 550
rect 0 31 50 469
<< mvndiff >>
rect 81 550 519 553
rect 81 494 519 500
rect 81 477 87 494
rect 513 477 519 494
rect 81 471 519 477
rect 79 469 521 471
rect -3 31 0 469
rect 50 463 521 469
rect 50 37 56 463
rect 73 415 521 463
rect 73 85 135 415
rect 465 85 521 415
rect 73 37 521 85
rect 50 31 521 37
rect 79 29 521 31
rect 81 23 519 29
rect 81 6 87 23
rect 513 6 519 23
rect 81 0 519 6
<< mvndiffc >>
rect 87 477 513 494
rect 56 37 73 463
rect 87 6 513 23
<< mvpsubdiff >>
rect 135 403 465 415
rect 135 97 147 403
rect 453 97 465 403
rect 135 85 465 97
rect 775 17 787 550
rect 1063 17 1075 550
rect 775 0 1075 17
<< mvpsubdiffcont >>
rect 147 97 453 403
rect 787 17 1063 550
<< poly >>
rect 0 542 81 550
rect 0 508 8 542
rect 42 508 81 542
rect 0 500 81 508
rect 519 542 600 550
rect 519 508 558 542
rect 592 508 600 542
rect 519 500 600 508
rect 0 469 50 500
rect 0 0 50 31
rect 550 0 600 500
<< polycont >>
rect 8 508 42 542
rect 558 508 592 542
<< locali >>
rect 0 542 50 550
rect 0 508 8 542
rect 42 508 50 542
rect 0 500 50 508
rect 550 542 600 550
rect 550 508 558 542
rect 592 508 600 542
rect 550 500 600 508
rect 79 477 87 494
rect 513 477 521 494
rect 73 471 527 477
rect 56 463 527 471
rect 73 415 527 463
rect 73 85 135 415
rect 465 85 527 415
rect 73 37 527 85
rect 56 29 527 37
rect 73 23 527 29
rect 79 6 87 23
rect 513 6 521 23
rect 775 17 787 550
rect 1063 17 1075 550
rect 775 0 1075 17
<< viali >>
rect 8 508 42 542
rect 558 508 592 542
rect 87 477 513 494
rect 56 37 73 463
rect 135 403 465 415
rect 135 97 147 403
rect 147 97 453 403
rect 453 97 465 403
rect 135 85 465 97
rect 87 6 513 23
rect 787 19 1063 550
<< metal1 >>
rect 0 542 50 550
rect 0 508 8 542
rect 42 508 50 542
rect 0 500 50 508
rect 550 542 600 550
rect 550 508 558 542
rect 592 508 600 542
rect 550 500 600 508
rect 81 494 519 497
rect 81 477 87 494
rect 513 477 519 494
rect 81 474 519 477
rect 76 469 524 474
rect 53 463 524 469
rect 53 37 56 463
rect 73 415 524 463
rect 73 85 135 415
rect 465 85 524 415
rect 73 37 524 85
rect 53 31 524 37
rect 76 26 524 31
rect 81 23 519 26
rect 81 6 87 23
rect 513 6 519 23
rect 81 3 519 6
rect 775 19 787 550
rect 1063 19 1075 550
rect 775 0 1075 19
<< via1 >>
rect 8 508 42 542
rect 558 508 592 542
rect 135 85 465 415
rect 875 38 975 138
<< metal2 >>
rect 0 542 775 550
rect 0 508 8 542
rect 42 508 558 542
rect 592 508 775 542
rect 0 500 775 508
rect 0 0 50 500
rect 125 415 475 425
rect 125 85 135 415
rect 465 85 475 415
rect 125 75 475 85
rect 550 0 775 500
rect 865 138 985 148
rect 865 38 875 138
rect 975 38 985 138
rect 865 28 985 38
<< via2 >>
rect 240 190 360 310
rect 875 38 975 138
<< metal3 >>
rect 0 510 226 550
tri 226 510 266 550 sw
tri 324 510 364 550 ne
rect 364 510 1075 550
rect 0 412 266 510
tri 266 412 364 510 sw
tri 364 412 462 510 ne
rect 462 412 1075 510
rect 0 324 364 412
tri 0 226 98 324 ne
rect 98 314 364 324
tri 364 314 462 412 sw
rect 98 310 1575 314
rect 98 226 240 310
tri 0 138 88 226 sw
tri 98 138 186 226 ne
rect 186 190 240 226
rect 360 190 1575 310
rect 186 138 1575 190
rect 0 58 88 138
tri 88 58 168 138 sw
tri 186 58 266 138 ne
rect 266 58 875 138
rect 0 0 168 58
tri 168 0 226 58 sw
tri 266 0 324 58 ne
rect 324 38 875 58
rect 975 38 1575 138
rect 324 0 1575 38
<< via3 >>
rect 240 190 360 310
rect 875 38 975 138
<< metal4 >>
rect 0 510 226 550
tri 226 510 266 550 sw
tri 324 510 364 550 ne
rect 364 510 1075 550
rect 0 412 266 510
tri 266 412 364 510 sw
tri 364 412 462 510 ne
rect 462 412 1075 510
rect 0 324 364 412
tri 0 226 98 324 ne
rect 98 314 364 324
tri 364 314 462 412 sw
rect 98 310 1575 314
rect 98 226 240 310
tri 0 138 88 226 sw
tri 98 138 186 226 ne
rect 186 190 240 226
rect 360 190 1575 310
rect 186 138 1575 190
rect 0 58 88 138
tri 88 58 168 138 sw
tri 186 58 266 138 ne
rect 266 58 875 138
rect 0 0 168 58
tri 168 0 226 58 sw
tri 266 0 324 58 ne
rect 324 38 875 58
rect 975 38 1575 138
rect 324 0 1575 38
<< via4 >>
rect 240 190 360 310
<< metal5 >>
rect 0 447 156 550
tri 156 447 259 550 sw
tri 394 447 497 550 ne
rect 497 447 1075 550
rect 0 394 259 447
tri 0 156 238 394 ne
rect 238 310 259 394
tri 259 310 396 447 sw
rect 238 190 240 310
rect 360 208 396 310
tri 396 208 498 310 sw
rect 360 190 1575 208
rect 238 156 1575 190
tri 0 0 156 156 sw
tri 238 0 394 156 ne
rect 394 0 1575 156
<< properties >>
string MASKHINTS_HVI 0 0 280 280 0 1920 280 2200
string MASKHINTS_HVNTM 2158 42 2214 1958
<< end >>
