magic
tech sky130A
timestamp 1693601174
<< checkpaint >>
rect -6555 -6605 25305 25255
<< dnwell >>
rect -3475 -3525 22225 22175
<< nwell >>
rect -5925 19825 24675 24625
rect -5925 -1175 -1125 19825
rect 19875 -1175 24675 19825
rect -5925 -5975 24675 -1175
<< pwell >>
rect -1125 18700 0 19825
rect 18700 18700 19875 19825
rect -1125 -1175 0 0
rect 18700 -1175 19875 0
<< mvnmos >>
rect 18700 18731 18750 19169
rect -469 -50 -31 0
rect 18781 -50 19219 0
rect 18700 -519 18750 -81
<< mvndiff >>
rect 18779 19169 19221 19171
rect -29 19163 0 19169
rect -29 18764 -23 19163
rect -64 18737 -23 18764
rect -6 18737 0 19163
rect -64 18731 0 18737
rect 18697 18731 18700 19169
rect 18750 19163 19221 19169
rect 18750 18737 18756 19163
rect 18773 19115 19221 19163
rect 18773 18785 18835 19115
rect 19165 18785 19221 19115
rect 18773 18737 19221 18785
rect 18750 18731 19221 18737
rect -64 18729 -31 18731
rect -469 18723 -31 18729
rect -469 18706 -463 18723
rect -37 18706 -31 18723
rect -469 18700 -31 18706
rect 18779 18729 19221 18731
rect 18781 18723 19219 18729
rect 18781 18706 18787 18723
rect 19213 18706 19219 18723
rect 18781 18700 19219 18706
rect -469 0 -31 3
rect 18781 0 19219 3
rect -469 -56 -31 -50
rect -469 -73 -463 -56
rect -37 -73 -31 -56
rect -469 -79 -31 -73
rect -471 -81 -29 -79
rect 18781 -56 19219 -50
rect 18781 -73 18787 -56
rect 19213 -73 19219 -56
rect 18781 -79 19219 -73
rect 18781 -81 18814 -79
rect -471 -87 0 -81
rect -471 -135 -23 -87
rect -471 -465 -415 -135
rect -85 -465 -23 -135
rect -471 -513 -23 -465
rect -6 -513 0 -87
rect -471 -519 0 -513
rect 18697 -519 18700 -81
rect 18750 -87 18814 -81
rect 18750 -513 18756 -87
rect 18773 -114 18814 -87
rect 18773 -513 18779 -114
rect 18750 -519 18779 -513
rect -471 -521 -29 -519
<< mvndiffc >>
rect -23 18737 -6 19163
rect 18756 18737 18773 19163
rect -463 18706 -37 18723
rect 18787 18706 19213 18723
rect -463 -73 -37 -56
rect 18787 -73 19213 -56
rect -23 -513 -6 -87
rect 18756 -513 18773 -87
<< mvpsubdiff >>
rect -1025 19713 0 19725
rect -1025 18717 -1013 19713
rect -19 19437 0 19713
rect -737 19425 0 19437
rect 18700 19713 19775 19725
rect 18700 19425 19487 19437
rect -737 18717 -725 19425
rect -1025 18700 -725 18717
rect 18835 19103 19165 19115
rect 18835 18797 18847 19103
rect 19153 18797 19165 19103
rect 18835 18785 19165 18797
rect 19475 18717 19487 19425
rect 19763 18717 19775 19713
rect 19475 18700 19775 18717
rect -1025 -1063 -1013 0
rect -737 -775 -725 0
rect -415 -147 -85 -135
rect -415 -453 -403 -147
rect -97 -453 -85 -147
rect -415 -465 -85 -453
rect 19475 -775 19487 0
rect -737 -787 0 -775
rect -17 -1063 0 -787
rect -1025 -1075 0 -1063
rect 18700 -787 19487 -775
rect 19763 -1063 19775 0
rect 18700 -1075 19775 -1063
<< mvnsubdiff >>
rect -5525 24213 24275 24225
rect -5525 -5563 -5513 24213
rect -1537 20225 20287 20237
rect -1537 -1575 -1525 20225
rect 20275 -1575 20287 20225
rect -1537 -1587 20287 -1575
rect 24263 -5563 24275 24213
rect -5525 -5575 24275 -5563
<< mvpsubdiffcont >>
rect -1013 19437 -19 19713
rect -1013 18717 -737 19437
rect 18700 19437 19763 19713
rect 18847 18797 19153 19103
rect 19487 18717 19763 19437
rect -1013 -787 -737 0
rect -403 -453 -97 -147
rect -1013 -1063 -17 -787
rect 19487 -787 19763 0
rect 18700 -1063 19763 -787
<< mvnsubdiffcont >>
rect -5513 20237 24263 24213
rect -5513 -1587 -1537 20237
rect 20287 -1587 24263 20237
rect -5513 -5563 24263 -1587
<< poly >>
rect -550 19242 0 19250
rect -550 19208 -542 19242
rect -508 19208 0 19242
rect -550 19200 0 19208
rect 18700 19242 19300 19250
rect 18700 19208 18708 19242
rect 18742 19208 19258 19242
rect 19292 19208 19300 19242
rect 18700 19200 19300 19208
rect -550 18700 -500 19200
rect 18700 19169 18750 19200
rect 18700 18700 18750 18731
rect 19250 18700 19300 19200
rect -550 -8 -469 0
rect -550 -42 -542 -8
rect -508 -42 -469 -8
rect -550 -50 -469 -42
rect -31 -50 0 0
rect 18700 -8 18781 0
rect 18700 -42 18708 -8
rect 18742 -42 18781 -8
rect 18700 -50 18781 -42
rect 19219 -8 19300 0
rect 19219 -42 19258 -8
rect 19292 -42 19300 -8
rect 19219 -50 19300 -42
rect -550 -550 -500 -50
rect 18700 -81 18750 -50
rect 18700 -550 18750 -519
rect 19250 -550 19300 -50
rect -550 -558 0 -550
rect -550 -592 -542 -558
rect -508 -592 0 -558
rect -550 -600 0 -592
rect 18700 -558 19300 -550
rect 18700 -592 18708 -558
rect 18742 -592 19258 -558
rect 19292 -592 19300 -558
rect 18700 -600 19300 -592
<< polycont >>
rect -542 19208 -508 19242
rect 18708 19208 18742 19242
rect 19258 19208 19292 19242
rect -542 -42 -508 -8
rect 18708 -42 18742 -8
rect 19258 -42 19292 -8
rect -542 -592 -508 -558
rect 18708 -592 18742 -558
rect 19258 -592 19292 -558
<< locali >>
rect -5525 24213 24275 24225
rect -5525 -5563 -5513 24213
rect -1537 20225 20287 20237
rect -1537 -1575 -1525 20225
rect -1025 19713 0 19725
rect -1025 18717 -1013 19713
rect -19 19437 0 19713
rect -737 19425 0 19437
rect 18700 19713 19775 19725
rect 18700 19425 19487 19437
rect -737 18717 -725 19425
rect -550 19242 -500 19250
rect -550 19208 -542 19242
rect -508 19208 -500 19242
rect -550 19200 -500 19208
rect 18700 19242 18750 19250
rect 18700 19208 18708 19242
rect 18742 19208 18750 19242
rect 18700 19200 18750 19208
rect 19250 19242 19300 19250
rect 19250 19208 19258 19242
rect 19292 19208 19300 19242
rect 19250 19200 19300 19208
rect 18773 19171 19227 19177
rect -23 19163 -6 19171
rect -64 18737 -23 18764
rect -64 18729 -6 18737
rect 18756 19163 19227 19171
rect 18773 19115 19227 19163
rect 18773 18785 18835 19115
rect 19165 18785 19227 19115
rect 18773 18737 19227 18785
rect 18756 18729 19227 18737
rect -64 18723 -29 18729
rect 18773 18723 19227 18729
rect -1025 18700 -725 18717
rect -471 18706 -463 18723
rect -37 18706 -29 18723
rect 18779 18706 18787 18723
rect 19213 18706 19221 18723
rect 19475 18717 19487 19425
rect 19763 18717 19775 19713
rect 19475 18700 19775 18717
rect -1025 -1063 -1013 0
rect -737 -775 -725 0
rect -550 -8 -500 0
rect -550 -42 -542 -8
rect -508 -42 -500 -8
rect -550 -50 -500 -42
rect 18700 -8 18750 0
rect 18700 -42 18708 -8
rect 18742 -42 18750 -8
rect 18700 -50 18750 -42
rect 19250 -8 19300 0
rect 19250 -42 19258 -8
rect 19292 -42 19300 -8
rect 19250 -50 19300 -42
rect -471 -73 -463 -56
rect -37 -73 -29 -56
rect 18779 -73 18787 -56
rect 19213 -73 19221 -56
rect -477 -79 -23 -73
rect 18779 -79 18814 -73
rect -477 -87 -6 -79
rect -477 -135 -23 -87
rect -477 -465 -415 -135
rect -85 -465 -23 -135
rect -477 -513 -23 -465
rect -477 -521 -6 -513
rect 18756 -87 18814 -79
rect 18773 -114 18814 -87
rect 18756 -521 18773 -513
rect -477 -527 -23 -521
rect -550 -558 -500 -550
rect -550 -592 -542 -558
rect -508 -592 -500 -558
rect -550 -600 -500 -592
rect 18700 -558 18750 -550
rect 18700 -592 18708 -558
rect 18742 -592 18750 -558
rect 18700 -600 18750 -592
rect 19250 -558 19300 -550
rect 19250 -592 19258 -558
rect 19292 -592 19300 -558
rect 19250 -600 19300 -592
rect 19475 -775 19487 0
rect -737 -787 0 -775
rect -17 -1063 0 -787
rect -1025 -1075 0 -1063
rect 18700 -787 19487 -775
rect 19763 -1063 19775 0
rect 18700 -1075 19775 -1063
rect 20275 -1575 20287 20225
rect -1537 -1587 20287 -1575
rect 24263 -5563 24275 24213
rect -5525 -5575 24275 -5563
<< viali >>
rect -5513 20237 24263 24213
rect -5513 -1587 -1537 20237
rect -1013 19437 -19 19713
rect -1013 18719 -737 19437
rect 18700 19437 19763 19713
rect -542 19208 -508 19242
rect 18708 19208 18742 19242
rect 19258 19208 19292 19242
rect -23 18737 -6 19163
rect 18756 18737 18773 19163
rect 18835 19103 19165 19115
rect 18835 18797 18847 19103
rect 18847 18797 19153 19103
rect 19153 18797 19165 19103
rect 18835 18785 19165 18797
rect -463 18706 -37 18723
rect 18787 18706 19213 18723
rect 19487 18719 19763 19437
rect -1013 -787 -737 0
rect -542 -42 -508 -8
rect 18708 -42 18742 -8
rect 19258 -42 19292 -8
rect -463 -73 -37 -56
rect 18787 -73 19213 -56
rect -415 -147 -85 -135
rect -415 -453 -403 -147
rect -403 -453 -97 -147
rect -97 -453 -85 -147
rect -415 -465 -85 -453
rect -23 -513 -6 -87
rect 18756 -513 18773 -87
rect -542 -592 -508 -558
rect 18708 -592 18742 -558
rect 19258 -592 19292 -558
rect -1013 -1063 -19 -787
rect 19487 -787 19763 0
rect 18700 -1063 19763 -787
rect 20287 -1587 24263 20237
rect -5513 -5563 24263 -1587
<< metal1 >>
rect -5525 24213 24275 24225
rect -5525 -5563 -5513 24213
rect -1537 20225 20287 20237
rect -1537 -1575 -1525 20225
rect -1025 19713 0 19725
rect -1025 18719 -1013 19713
rect -19 19437 0 19713
rect -737 19425 0 19437
rect 18700 19713 19775 19725
rect 18700 19425 19487 19437
rect -737 18719 -725 19425
rect -550 19242 -500 19250
rect -550 19208 -542 19242
rect -508 19208 -500 19242
rect -550 19200 -500 19208
rect 18700 19242 18750 19250
rect 18700 19208 18708 19242
rect 18742 19208 18750 19242
rect 18700 19200 18750 19208
rect 19250 19242 19300 19250
rect 19250 19208 19258 19242
rect 19292 19208 19300 19242
rect 19250 19200 19300 19208
rect -474 19169 -26 19174
rect 18776 19169 19224 19174
rect -474 19163 -3 19169
rect -474 19115 -23 19163
rect -474 18785 -415 19115
rect -85 18785 -23 19115
rect -474 18737 -23 18785
rect -6 18737 -3 19163
rect -474 18731 -3 18737
rect 18753 19163 19224 19169
rect 18753 18737 18756 19163
rect 18773 19115 19224 19163
rect 18773 18785 18835 19115
rect 19165 18785 19224 19115
rect 18773 18737 19224 18785
rect 18753 18731 19224 18737
rect -474 18726 -26 18731
rect 18776 18726 19224 18731
rect -1025 18700 -725 18719
rect -469 18723 -31 18726
rect -469 18706 -463 18723
rect -37 18706 -31 18723
rect -469 18703 -31 18706
rect 18781 18723 19219 18726
rect 18781 18706 18787 18723
rect 19213 18706 19219 18723
rect 18781 18703 19219 18706
rect 19475 18719 19487 19425
rect 19763 18719 19775 19713
rect 19475 18700 19775 18719
rect -1025 -1063 -1013 0
rect -737 -775 -725 0
rect -550 -8 -500 0
rect -550 -42 -542 -8
rect -508 -42 -500 -8
rect -550 -50 -500 -42
rect 18700 -8 18750 0
rect 18700 -42 18708 -8
rect 18742 -42 18750 -8
rect 18700 -50 18750 -42
rect 19250 -8 19300 0
rect 19250 -42 19258 -8
rect 19292 -42 19300 -8
rect 19250 -50 19300 -42
rect -469 -56 -31 -53
rect -469 -73 -463 -56
rect -37 -73 -31 -56
rect -469 -76 -31 -73
rect 18781 -56 19219 -53
rect 18781 -73 18787 -56
rect 19213 -73 19219 -56
rect 18781 -76 19219 -73
rect -474 -81 -26 -76
rect 18776 -81 19224 -76
rect -474 -87 -3 -81
rect -474 -135 -23 -87
rect -474 -465 -415 -135
rect -85 -465 -23 -135
rect -474 -513 -23 -465
rect -6 -513 -3 -87
rect -474 -519 -3 -513
rect 18753 -87 19224 -81
rect 18753 -513 18756 -87
rect 18773 -135 19224 -87
rect 18773 -465 18835 -135
rect 19165 -465 19224 -135
rect 18773 -513 19224 -465
rect 18753 -519 19224 -513
rect -474 -524 -26 -519
rect 18776 -524 19224 -519
rect -550 -558 -500 -550
rect -550 -592 -542 -558
rect -508 -592 -500 -558
rect -550 -600 -500 -592
rect 18700 -558 18750 -550
rect 18700 -592 18708 -558
rect 18742 -592 18750 -558
rect 18700 -600 18750 -592
rect 19250 -558 19300 -550
rect 19250 -592 19258 -558
rect 19292 -592 19300 -558
rect 19250 -600 19300 -592
rect 19475 -775 19487 0
rect -737 -787 0 -775
rect -19 -1063 0 -787
rect -1025 -1075 0 -1063
rect 18700 -787 19487 -775
rect 19763 -1063 19775 0
rect 18700 -1075 19775 -1063
rect 20275 -1575 20287 20225
rect -1537 -1587 20287 -1575
rect 24263 -5563 24275 24213
rect -5525 -5575 24275 -5563
<< via1 >>
rect -5513 20237 24263 24213
rect -5513 1117 -1537 20225
rect 18788 19525 18888 19625
rect -542 19208 -508 19242
rect 18708 19208 18742 19242
rect 19258 19208 19292 19242
rect -415 18785 -85 19115
rect 18835 18785 19165 19115
rect 19575 18738 19675 18838
rect -925 -188 -825 -88
rect -542 -42 -508 -8
rect 18708 -42 18742 -8
rect 19258 -42 19292 -8
rect -415 -465 -85 -135
rect 18835 -465 19165 -135
rect -542 -592 -508 -558
rect 18708 -592 18742 -558
rect 19258 -592 19292 -558
rect -138 -975 -38 -875
rect 20287 -1587 24263 20237
rect -495 -5563 24263 -1587
<< metal2 >>
rect -5525 24213 24275 24225
rect -5525 20237 -5513 24213
rect -5525 20225 20287 20237
rect -5525 1117 -5513 20225
rect -1537 1117 -1525 20225
rect 18778 19625 18898 19635
rect 18778 19525 18788 19625
rect 18888 19525 18898 19625
rect 18778 19515 18898 19525
rect -725 19242 0 19425
rect -725 19208 -542 19242
rect -508 19208 0 19242
rect -725 19200 0 19208
rect 18700 19242 19475 19425
rect 18700 19208 18708 19242
rect 18742 19208 19258 19242
rect 19292 19208 19475 19242
rect 18700 19200 19475 19208
rect -725 18700 -500 19200
rect -425 19115 -75 19125
rect -425 18785 -415 19115
rect -85 18785 -75 19115
rect -425 18775 -75 18785
rect 18700 18700 18750 19200
rect 18825 19115 19175 19125
rect 18825 18785 18835 19115
rect 19165 18785 19175 19115
rect 18825 18775 19175 18785
rect 19250 18700 19475 19200
rect 19565 18838 19685 18848
rect 19565 18738 19575 18838
rect 19675 18738 19685 18838
rect 19565 18728 19685 18738
rect -725 -8 0 0
rect -725 -42 -542 -8
rect -508 -42 0 -8
rect -725 -50 0 -42
rect 18700 -8 19475 0
rect 18700 -42 18708 -8
rect 18742 -42 19258 -8
rect 19292 -42 19475 -8
rect 18700 -50 19475 -42
rect -935 -88 -815 -78
rect -935 -188 -925 -88
rect -825 -188 -815 -88
rect -935 -198 -815 -188
rect -725 -550 -500 -50
rect -425 -135 -75 -125
rect -425 -465 -415 -135
rect -85 -465 -75 -135
rect -425 -475 -75 -465
rect 18700 -550 18750 -50
rect 18825 -135 19175 -125
rect 18825 -465 18835 -135
rect 19165 -465 19175 -135
rect 18825 -475 19175 -465
rect 19250 -550 19475 -50
rect -725 -558 0 -550
rect -725 -592 -542 -558
rect -508 -592 0 -558
rect -725 -775 0 -592
rect 18700 -558 19475 -550
rect 18700 -592 18708 -558
rect 18742 -592 19258 -558
rect 19292 -592 19475 -558
rect 18700 -775 19475 -592
rect -148 -875 -28 -865
rect -148 -975 -138 -875
rect -38 -975 -28 -875
rect -148 -985 -28 -975
rect 20275 -1575 20287 20225
rect -507 -1587 20287 -1575
rect -507 -5563 -495 -1587
rect 24263 -5563 24275 24213
rect -507 -5575 24275 -5563
<< via2 >>
rect 18788 19525 18888 19625
rect -310 18890 -190 19010
rect 18940 18890 19060 19010
rect 19575 18738 19675 18838
rect -925 -188 -825 -88
rect -310 -360 -190 -240
rect 18940 -360 19060 -240
rect -138 -975 -38 -875
<< metal3 >>
rect -2525 20225 19275 21225
rect -2525 19338 -1525 20225
rect -638 19338 -186 20225
rect -2525 19014 -186 19338
rect -88 19112 0 19725
tri -186 19014 -88 19112 sw
tri -88 19024 0 19112 ne
rect 18700 19625 19064 19725
rect 18700 19525 18788 19625
rect 18888 19525 19064 19625
rect 18700 19024 19064 19525
tri 18700 19014 18710 19024 ne
rect 18710 19014 19064 19024
tri 19064 19014 19162 19112 sw
rect 20275 19014 21275 19225
rect -2525 19010 -88 19014
rect -2525 18890 -310 19010
rect -190 18926 -88 19010
tri -88 18926 0 19014 sw
tri 18710 18926 18798 19014 ne
rect 18798 19010 21275 19014
rect 18798 18926 18940 19010
rect -190 18890 0 18926
rect -2525 18886 0 18890
rect -2525 -575 -1525 18886
tri -412 18788 -314 18886 ne
rect -314 18788 0 18886
rect -1025 18700 -412 18788
tri -412 18700 -324 18788 sw
tri -314 18700 -226 18788 ne
rect -226 18700 0 18788
tri 18700 18838 18788 18926 sw
tri 18798 18838 18886 18926 ne
rect 18886 18890 18940 18926
rect 19060 18890 21275 19010
rect 18886 18838 21275 18890
rect 18700 18758 18788 18838
tri 18788 18758 18868 18838 sw
tri 18886 18758 18966 18838 ne
rect 18966 18758 19575 18838
rect 18700 18700 18868 18758
tri 18868 18700 18926 18758 sw
tri 18966 18700 19024 18758 ne
rect 19024 18738 19575 18758
rect 19675 18738 21275 18838
rect 19024 18700 21275 18738
rect 20275 0 21275 18700
rect -1025 -40 -324 0
tri -324 -40 -284 0 sw
tri -226 -40 -186 0 ne
rect -186 -40 0 0
rect -1025 -88 -284 -40
rect -1025 -188 -925 -88
rect -825 -138 -284 -88
tri -284 -138 -186 -40 sw
tri -186 -138 -88 -40 ne
rect -88 -138 0 -40
rect -825 -188 -186 -138
rect -1025 -236 -186 -188
tri -186 -236 -88 -138 sw
tri -88 -226 0 -138 ne
rect 18700 -40 18926 0
tri 18926 -40 18966 0 sw
tri 19024 -40 19064 0 ne
rect 19064 -40 21275 0
rect 18700 -138 18966 -40
tri 18966 -138 19064 -40 sw
tri 19064 -138 19162 -40 ne
rect 19162 -138 21275 -40
rect 18700 -226 19064 -138
tri 18700 -236 18710 -226 ne
rect 18710 -236 19064 -226
tri 19064 -236 19162 -138 sw
rect -1025 -240 -88 -236
rect -1025 -360 -310 -240
rect -190 -324 -88 -240
tri -88 -324 0 -236 sw
tri 18710 -324 18798 -236 ne
rect 18798 -240 19775 -236
rect 18798 -324 18940 -240
rect -190 -360 0 -324
rect -1025 -364 0 -360
tri -412 -462 -314 -364 ne
rect -314 -875 0 -364
rect -314 -975 -138 -875
rect -38 -975 0 -875
rect -314 -1575 0 -975
tri 18700 -364 18740 -324 sw
tri 18798 -364 18838 -324 ne
rect 18838 -360 18940 -324
rect 19060 -360 19775 -240
rect 18838 -364 19775 -360
rect 18700 -462 18740 -364
tri 18740 -462 18838 -364 sw
tri 18838 -462 18936 -364 ne
rect 18700 -1575 18838 -462
rect 18936 -688 19775 -364
rect 18936 -1075 19388 -688
rect 20275 -1575 21275 -138
rect -525 -2575 21275 -1575
<< via3 >>
rect 18788 19525 18888 19625
rect -310 18890 -190 19010
rect 18940 18890 19060 19010
rect 19575 18738 19675 18838
rect -925 -188 -825 -88
rect -310 -360 -190 -240
rect -138 -975 -38 -875
rect 18940 -360 19060 -240
<< metal4 >>
rect -2525 20225 19275 21225
rect -2525 19338 -1525 20225
rect -638 19338 -186 20225
rect -2525 19014 -186 19338
rect -88 19112 0 19725
tri -186 19014 -88 19112 sw
tri -88 19024 0 19112 ne
rect 18700 19625 19064 19725
rect 18700 19525 18788 19625
rect 18888 19525 19064 19625
rect 18700 19024 19064 19525
tri 18700 19014 18710 19024 ne
rect 18710 19014 19064 19024
tri 19064 19014 19162 19112 sw
rect 20275 19014 21275 19225
rect -2525 19010 -88 19014
rect -2525 18890 -310 19010
rect -190 18926 -88 19010
tri -88 18926 0 19014 sw
tri 18710 18926 18798 19014 ne
rect 18798 19010 21275 19014
rect 18798 18926 18940 19010
rect -190 18890 0 18926
rect -2525 18886 0 18890
rect -2525 -575 -1525 18886
tri -412 18788 -314 18886 ne
rect -314 18788 0 18886
rect -1025 18700 -412 18788
tri -412 18700 -324 18788 sw
tri -314 18700 -226 18788 ne
rect -226 18700 0 18788
tri 18700 18838 18788 18926 sw
tri 18798 18838 18886 18926 ne
rect 18886 18890 18940 18926
rect 19060 18890 21275 19010
rect 18886 18838 21275 18890
rect 18700 18758 18788 18838
tri 18788 18758 18868 18838 sw
tri 18886 18758 18966 18838 ne
rect 18966 18758 19575 18838
rect 18700 18700 18868 18758
tri 18868 18700 18926 18758 sw
tri 18966 18700 19024 18758 ne
rect 19024 18738 19575 18758
rect 19675 18738 21275 18838
rect 19024 18700 21275 18738
rect 20275 0 21275 18700
rect -1025 -40 -324 0
tri -324 -40 -284 0 sw
tri -226 -40 -186 0 ne
rect -186 -40 0 0
rect -1025 -88 -284 -40
rect -1025 -188 -925 -88
rect -825 -138 -284 -88
tri -284 -138 -186 -40 sw
tri -186 -138 -88 -40 ne
rect -88 -138 0 -40
rect -825 -188 -186 -138
rect -1025 -236 -186 -188
tri -186 -236 -88 -138 sw
tri -88 -226 0 -138 ne
rect 18700 -40 18926 0
tri 18926 -40 18966 0 sw
tri 19024 -40 19064 0 ne
rect 19064 -40 21275 0
rect 18700 -138 18966 -40
tri 18966 -138 19064 -40 sw
tri 19064 -138 19162 -40 ne
rect 19162 -138 21275 -40
rect 18700 -226 19064 -138
tri 18700 -236 18710 -226 ne
rect 18710 -236 19064 -226
tri 19064 -236 19162 -138 sw
rect -1025 -240 -88 -236
rect -1025 -360 -310 -240
rect -190 -324 -88 -240
tri -88 -324 0 -236 sw
tri 18710 -324 18798 -236 ne
rect 18798 -240 19775 -236
rect 18798 -324 18940 -240
rect -190 -360 0 -324
rect -1025 -364 0 -360
tri -412 -462 -314 -364 ne
rect -314 -875 0 -364
rect -314 -975 -138 -875
rect -38 -975 0 -875
rect -314 -1575 0 -975
tri 18700 -364 18740 -324 sw
tri 18798 -364 18838 -324 ne
rect 18838 -360 18940 -324
rect 19060 -360 19775 -240
rect 18838 -364 19775 -360
rect 18700 -462 18740 -364
tri 18740 -462 18838 -364 sw
tri 18838 -462 18936 -364 ne
rect 18700 -1575 18838 -462
rect 18936 -688 19775 -364
rect 18936 -1075 19388 -688
rect 20275 -1575 21275 -138
rect -525 -2575 21275 -1575
<< via4 >>
rect -310 18890 -190 19010
rect 18940 18890 19060 19010
rect -310 -360 -190 -240
rect 18940 -360 19060 -240
<< metal5 >>
rect -2525 20225 19275 21225
rect -2525 19303 -1525 20225
rect -603 19303 -292 20225
rect -2525 19010 -292 19303
tri -292 19010 -154 19148 sw
rect -53 19147 0 19725
tri -53 19094 0 19147 ne
rect 18700 19094 18958 19725
tri 18700 19010 18784 19094 ne
rect 18784 19010 18958 19094
tri 18958 19010 19096 19148 sw
rect -2525 18992 -310 19010
rect -2525 -575 -1525 18992
tri -448 18890 -346 18992 ne
rect -346 18890 -310 18992
rect -190 18890 -154 19010
tri -346 18753 -209 18890 ne
rect -209 18856 -154 18890
tri -154 18856 0 19010 sw
tri 18784 18856 18938 19010 ne
rect 18938 18890 18940 19010
rect 19060 18908 19096 19010
tri 19096 18908 19198 19010 sw
rect 20275 18908 21275 19225
rect 19060 18890 21275 18908
rect 18938 18856 21275 18890
rect -209 18753 0 18856
rect -1025 18700 -447 18753
tri -447 18700 -394 18753 sw
tri -209 18700 -156 18753 ne
rect -156 18700 0 18753
tri 18700 18700 18856 18856 sw
tri 18938 18700 19094 18856 ne
rect 19094 18700 21275 18856
rect 20275 0 21275 18700
rect -1025 -103 -394 0
tri -394 -103 -291 0 sw
tri -156 -103 -53 0 ne
rect -53 -103 0 0
rect -1025 -240 -291 -103
tri -291 -240 -154 -103 sw
tri -53 -156 0 -103 ne
rect 18700 -103 18856 0
tri 18856 -103 18959 0 sw
tri 19094 -103 19197 0 ne
rect 19197 -103 21275 0
rect 18700 -156 18959 -103
tri 18700 -240 18784 -156 ne
rect 18784 -240 18959 -156
tri 18959 -240 19096 -103 sw
rect -1025 -258 -310 -240
tri -448 -360 -346 -258 ne
rect -346 -360 -310 -258
rect -190 -360 -154 -240
tri -346 -498 -208 -360 ne
rect -208 -394 -154 -360
tri -154 -394 0 -240 sw
tri 18784 -394 18938 -240 ne
rect 18938 -360 18940 -240
rect 19060 -342 19096 -240
tri 19096 -342 19198 -240 sw
rect 19060 -360 19775 -342
rect 18938 -394 19775 -360
rect -208 -1575 0 -394
tri 18700 -497 18803 -394 sw
rect 18700 -1575 18803 -497
tri 18938 -498 19042 -394 ne
rect 19042 -653 19775 -394
rect 19042 -1075 19353 -653
rect 20275 -1575 21275 -103
rect -525 -2575 21275 -1575
use nmos_drain_frame_lt  nmos_drain_frame_lt_0 waffle_cells
timestamp 1675431365
transform 1 0 -550 0 1 0
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_1
timestamp 1675431365
transform 0 -1 1100 -1 0 19250
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_2
timestamp 1675431365
transform 1 0 -550 0 1 1100
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_3
timestamp 1675431365
transform 0 -1 2200 -1 0 19250
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_4
timestamp 1675431365
transform 1 0 -550 0 1 2200
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_5
timestamp 1675431365
transform 0 -1 3300 -1 0 19250
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_6
timestamp 1675431365
transform 1 0 -550 0 1 3300
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_7
timestamp 1675431365
transform 0 -1 4400 -1 0 19250
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_8
timestamp 1675431365
transform 1 0 -550 0 1 4400
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_9
timestamp 1675431365
transform 0 -1 5500 -1 0 19250
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_10
timestamp 1675431365
transform 1 0 -550 0 1 5500
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_11
timestamp 1675431365
transform 0 -1 6600 -1 0 19250
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_12
timestamp 1675431365
transform 1 0 -550 0 1 6600
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_13
timestamp 1675431365
transform 0 -1 7700 -1 0 19250
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_14
timestamp 1675431365
transform 1 0 -550 0 1 7700
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_15
timestamp 1675431365
transform 0 -1 8800 -1 0 19250
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_16
timestamp 1675431365
transform 1 0 -550 0 1 8800
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_17
timestamp 1675431365
transform 0 -1 9900 -1 0 19250
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_18
timestamp 1675431365
transform 1 0 -550 0 1 9900
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_19
timestamp 1675431365
transform 0 -1 11000 -1 0 19250
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_20
timestamp 1675431365
transform 1 0 -550 0 1 11000
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_21
timestamp 1675431365
transform 0 -1 12100 -1 0 19250
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_22
timestamp 1675431365
transform 1 0 -550 0 1 12100
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_23
timestamp 1675431365
transform 0 -1 13200 -1 0 19250
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_24
timestamp 1675431365
transform 1 0 -550 0 1 13200
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_25
timestamp 1675431365
transform 0 -1 14300 -1 0 19250
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_26
timestamp 1675431365
transform 1 0 -550 0 1 14300
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_27
timestamp 1675431365
transform 0 -1 15400 -1 0 19250
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_28
timestamp 1675431365
transform 1 0 -550 0 1 15400
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_29
timestamp 1675431365
transform 0 -1 16500 -1 0 19250
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_30
timestamp 1675431365
transform 1 0 -550 0 1 16500
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_31
timestamp 1675431365
transform 0 -1 17600 -1 0 19250
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_32
timestamp 1675431365
transform 1 0 -550 0 1 17600
box -975 -113 663 663
use nmos_drain_frame_lt  nmos_drain_frame_lt_33
timestamp 1675431365
transform 0 -1 18700 -1 0 19250
box -975 -113 663 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_0 waffle_cells
timestamp 1675431051
transform 0 -1 550 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_1
timestamp 1675431051
transform 1 0 18700 0 1 550
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_2
timestamp 1675431051
transform 0 -1 1650 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_3
timestamp 1675431051
transform 1 0 18700 0 1 1650
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_4
timestamp 1675431051
transform 0 -1 2750 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_5
timestamp 1675431051
transform 1 0 18700 0 1 2750
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_6
timestamp 1675431051
transform 0 -1 3850 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_7
timestamp 1675431051
transform 1 0 18700 0 1 3850
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_8
timestamp 1675431051
transform 0 -1 4950 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_9
timestamp 1675431051
transform 1 0 18700 0 1 4950
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_10
timestamp 1675431051
transform 0 -1 6050 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_11
timestamp 1675431051
transform 1 0 18700 0 1 6050
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_12
timestamp 1675431051
transform 0 -1 7150 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_13
timestamp 1675431051
transform 1 0 18700 0 1 7150
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_14
timestamp 1675431051
transform 0 -1 8250 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_15
timestamp 1675431051
transform 1 0 18700 0 1 8250
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_16
timestamp 1675431051
transform 0 -1 9350 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_17
timestamp 1675431051
transform 1 0 18700 0 1 9350
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_18
timestamp 1675431051
transform 0 -1 10450 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_19
timestamp 1675431051
transform 1 0 18700 0 1 10450
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_20
timestamp 1675431051
transform 0 -1 11550 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_21
timestamp 1675431051
transform 1 0 18700 0 1 11550
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_22
timestamp 1675431051
transform 0 -1 12650 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_23
timestamp 1675431051
transform 1 0 18700 0 1 12650
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_24
timestamp 1675431051
transform 0 -1 13750 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_25
timestamp 1675431051
transform 1 0 18700 0 1 13750
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_26
timestamp 1675431051
transform 0 -1 14850 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_27
timestamp 1675431051
transform 1 0 18700 0 1 14850
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_28
timestamp 1675431051
transform 0 -1 15950 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_29
timestamp 1675431051
transform 1 0 18700 0 1 15950
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_30
timestamp 1675431051
transform 0 -1 17050 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_31
timestamp 1675431051
transform 1 0 18700 0 1 17050
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_32
timestamp 1675431051
transform 0 -1 18150 -1 0 0
box -113 -113 1575 663
use nmos_drain_frame_rb  nmos_drain_frame_rb_33
timestamp 1675431051
transform 1 0 18700 0 1 18150
box -113 -113 1575 663
use nmos_drain_in  nmos_drain_in_0 waffle_cells
timestamp 1675431861
transform 1 0 0 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_1
timestamp 1675431861
transform 1 0 0 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_2
timestamp 1675431861
transform 1 0 0 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_3
timestamp 1675431861
transform 1 0 0 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_4
timestamp 1675431861
transform 1 0 0 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_5
timestamp 1675431861
transform 1 0 0 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_6
timestamp 1675431861
transform 1 0 0 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_7
timestamp 1675431861
transform 1 0 0 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_8
timestamp 1675431861
transform 1 0 0 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_9
timestamp 1675431861
transform 1 0 0 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_10
timestamp 1675431861
transform 1 0 0 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_11
timestamp 1675431861
transform 1 0 0 0 1 12650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_12
timestamp 1675431861
transform 1 0 0 0 1 13750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_13
timestamp 1675431861
transform 1 0 0 0 1 14850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_14
timestamp 1675431861
transform 1 0 0 0 1 15950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_15
timestamp 1675431861
transform 1 0 0 0 1 17050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_16
timestamp 1675431861
transform 1 0 0 0 1 18150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_17
timestamp 1675431861
transform 1 0 550 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_18
timestamp 1675431861
transform 1 0 550 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_19
timestamp 1675431861
transform 1 0 550 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_20
timestamp 1675431861
transform 1 0 550 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_21
timestamp 1675431861
transform 1 0 550 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_22
timestamp 1675431861
transform 1 0 550 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_23
timestamp 1675431861
transform 1 0 550 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_24
timestamp 1675431861
transform 1 0 550 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_25
timestamp 1675431861
transform 1 0 550 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_26
timestamp 1675431861
transform 1 0 550 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_27
timestamp 1675431861
transform 1 0 550 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_28
timestamp 1675431861
transform 1 0 550 0 1 12100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_29
timestamp 1675431861
transform 1 0 550 0 1 13200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_30
timestamp 1675431861
transform 1 0 550 0 1 14300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_31
timestamp 1675431861
transform 1 0 550 0 1 15400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_32
timestamp 1675431861
transform 1 0 550 0 1 16500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_33
timestamp 1675431861
transform 1 0 550 0 1 17600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_34
timestamp 1675431861
transform 1 0 1100 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_35
timestamp 1675431861
transform 1 0 1100 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_36
timestamp 1675431861
transform 1 0 1100 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_37
timestamp 1675431861
transform 1 0 1100 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_38
timestamp 1675431861
transform 1 0 1100 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_39
timestamp 1675431861
transform 1 0 1100 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_40
timestamp 1675431861
transform 1 0 1100 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_41
timestamp 1675431861
transform 1 0 1100 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_42
timestamp 1675431861
transform 1 0 1100 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_43
timestamp 1675431861
transform 1 0 1100 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_44
timestamp 1675431861
transform 1 0 1100 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_45
timestamp 1675431861
transform 1 0 1100 0 1 12650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_46
timestamp 1675431861
transform 1 0 1100 0 1 13750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_47
timestamp 1675431861
transform 1 0 1100 0 1 14850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_48
timestamp 1675431861
transform 1 0 1100 0 1 15950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_49
timestamp 1675431861
transform 1 0 1100 0 1 17050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_50
timestamp 1675431861
transform 1 0 1100 0 1 18150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_51
timestamp 1675431861
transform 1 0 1650 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_52
timestamp 1675431861
transform 1 0 1650 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_53
timestamp 1675431861
transform 1 0 1650 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_54
timestamp 1675431861
transform 1 0 1650 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_55
timestamp 1675431861
transform 1 0 1650 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_56
timestamp 1675431861
transform 1 0 1650 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_57
timestamp 1675431861
transform 1 0 1650 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_58
timestamp 1675431861
transform 1 0 1650 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_59
timestamp 1675431861
transform 1 0 1650 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_60
timestamp 1675431861
transform 1 0 1650 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_61
timestamp 1675431861
transform 1 0 1650 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_62
timestamp 1675431861
transform 1 0 1650 0 1 12100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_63
timestamp 1675431861
transform 1 0 1650 0 1 13200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_64
timestamp 1675431861
transform 1 0 1650 0 1 14300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_65
timestamp 1675431861
transform 1 0 1650 0 1 15400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_66
timestamp 1675431861
transform 1 0 1650 0 1 16500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_67
timestamp 1675431861
transform 1 0 1650 0 1 17600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_68
timestamp 1675431861
transform 1 0 2200 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_69
timestamp 1675431861
transform 1 0 2200 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_70
timestamp 1675431861
transform 1 0 2200 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_71
timestamp 1675431861
transform 1 0 2200 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_72
timestamp 1675431861
transform 1 0 2200 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_73
timestamp 1675431861
transform 1 0 2200 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_74
timestamp 1675431861
transform 1 0 2200 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_75
timestamp 1675431861
transform 1 0 2200 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_76
timestamp 1675431861
transform 1 0 2200 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_77
timestamp 1675431861
transform 1 0 2200 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_78
timestamp 1675431861
transform 1 0 2200 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_79
timestamp 1675431861
transform 1 0 2200 0 1 12650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_80
timestamp 1675431861
transform 1 0 2200 0 1 13750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_81
timestamp 1675431861
transform 1 0 2200 0 1 14850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_82
timestamp 1675431861
transform 1 0 2200 0 1 15950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_83
timestamp 1675431861
transform 1 0 2200 0 1 17050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_84
timestamp 1675431861
transform 1 0 2200 0 1 18150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_85
timestamp 1675431861
transform 1 0 2750 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_86
timestamp 1675431861
transform 1 0 2750 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_87
timestamp 1675431861
transform 1 0 2750 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_88
timestamp 1675431861
transform 1 0 2750 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_89
timestamp 1675431861
transform 1 0 2750 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_90
timestamp 1675431861
transform 1 0 2750 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_91
timestamp 1675431861
transform 1 0 2750 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_92
timestamp 1675431861
transform 1 0 2750 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_93
timestamp 1675431861
transform 1 0 2750 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_94
timestamp 1675431861
transform 1 0 2750 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_95
timestamp 1675431861
transform 1 0 2750 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_96
timestamp 1675431861
transform 1 0 2750 0 1 12100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_97
timestamp 1675431861
transform 1 0 2750 0 1 13200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_98
timestamp 1675431861
transform 1 0 2750 0 1 14300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_99
timestamp 1675431861
transform 1 0 2750 0 1 15400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_100
timestamp 1675431861
transform 1 0 2750 0 1 16500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_101
timestamp 1675431861
transform 1 0 2750 0 1 17600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_102
timestamp 1675431861
transform 1 0 3300 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_103
timestamp 1675431861
transform 1 0 3300 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_104
timestamp 1675431861
transform 1 0 3300 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_105
timestamp 1675431861
transform 1 0 3300 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_106
timestamp 1675431861
transform 1 0 3300 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_107
timestamp 1675431861
transform 1 0 3300 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_108
timestamp 1675431861
transform 1 0 3300 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_109
timestamp 1675431861
transform 1 0 3300 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_110
timestamp 1675431861
transform 1 0 3300 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_111
timestamp 1675431861
transform 1 0 3300 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_112
timestamp 1675431861
transform 1 0 3300 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_113
timestamp 1675431861
transform 1 0 3300 0 1 12650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_114
timestamp 1675431861
transform 1 0 3300 0 1 13750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_115
timestamp 1675431861
transform 1 0 3300 0 1 14850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_116
timestamp 1675431861
transform 1 0 3300 0 1 15950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_117
timestamp 1675431861
transform 1 0 3300 0 1 17050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_118
timestamp 1675431861
transform 1 0 3300 0 1 18150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_119
timestamp 1675431861
transform 1 0 3850 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_120
timestamp 1675431861
transform 1 0 3850 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_121
timestamp 1675431861
transform 1 0 3850 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_122
timestamp 1675431861
transform 1 0 3850 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_123
timestamp 1675431861
transform 1 0 3850 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_124
timestamp 1675431861
transform 1 0 3850 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_125
timestamp 1675431861
transform 1 0 3850 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_126
timestamp 1675431861
transform 1 0 3850 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_127
timestamp 1675431861
transform 1 0 3850 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_128
timestamp 1675431861
transform 1 0 3850 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_129
timestamp 1675431861
transform 1 0 3850 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_130
timestamp 1675431861
transform 1 0 3850 0 1 12100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_131
timestamp 1675431861
transform 1 0 3850 0 1 13200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_132
timestamp 1675431861
transform 1 0 3850 0 1 14300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_133
timestamp 1675431861
transform 1 0 3850 0 1 15400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_134
timestamp 1675431861
transform 1 0 3850 0 1 16500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_135
timestamp 1675431861
transform 1 0 3850 0 1 17600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_136
timestamp 1675431861
transform 1 0 4400 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_137
timestamp 1675431861
transform 1 0 4400 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_138
timestamp 1675431861
transform 1 0 4400 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_139
timestamp 1675431861
transform 1 0 4400 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_140
timestamp 1675431861
transform 1 0 4400 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_141
timestamp 1675431861
transform 1 0 4400 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_142
timestamp 1675431861
transform 1 0 4400 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_143
timestamp 1675431861
transform 1 0 4400 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_144
timestamp 1675431861
transform 1 0 4400 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_145
timestamp 1675431861
transform 1 0 4400 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_146
timestamp 1675431861
transform 1 0 4400 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_147
timestamp 1675431861
transform 1 0 4400 0 1 12650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_148
timestamp 1675431861
transform 1 0 4400 0 1 13750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_149
timestamp 1675431861
transform 1 0 4400 0 1 14850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_150
timestamp 1675431861
transform 1 0 4400 0 1 15950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_151
timestamp 1675431861
transform 1 0 4400 0 1 17050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_152
timestamp 1675431861
transform 1 0 4400 0 1 18150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_153
timestamp 1675431861
transform 1 0 4950 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_154
timestamp 1675431861
transform 1 0 4950 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_155
timestamp 1675431861
transform 1 0 4950 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_156
timestamp 1675431861
transform 1 0 4950 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_157
timestamp 1675431861
transform 1 0 4950 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_158
timestamp 1675431861
transform 1 0 4950 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_159
timestamp 1675431861
transform 1 0 4950 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_160
timestamp 1675431861
transform 1 0 4950 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_161
timestamp 1675431861
transform 1 0 4950 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_162
timestamp 1675431861
transform 1 0 4950 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_163
timestamp 1675431861
transform 1 0 4950 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_164
timestamp 1675431861
transform 1 0 4950 0 1 12100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_165
timestamp 1675431861
transform 1 0 4950 0 1 13200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_166
timestamp 1675431861
transform 1 0 4950 0 1 14300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_167
timestamp 1675431861
transform 1 0 4950 0 1 15400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_168
timestamp 1675431861
transform 1 0 4950 0 1 16500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_169
timestamp 1675431861
transform 1 0 4950 0 1 17600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_170
timestamp 1675431861
transform 1 0 5500 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_171
timestamp 1675431861
transform 1 0 5500 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_172
timestamp 1675431861
transform 1 0 5500 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_173
timestamp 1675431861
transform 1 0 5500 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_174
timestamp 1675431861
transform 1 0 5500 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_175
timestamp 1675431861
transform 1 0 5500 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_176
timestamp 1675431861
transform 1 0 5500 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_177
timestamp 1675431861
transform 1 0 5500 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_178
timestamp 1675431861
transform 1 0 5500 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_179
timestamp 1675431861
transform 1 0 5500 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_180
timestamp 1675431861
transform 1 0 5500 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_181
timestamp 1675431861
transform 1 0 5500 0 1 12650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_182
timestamp 1675431861
transform 1 0 5500 0 1 13750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_183
timestamp 1675431861
transform 1 0 5500 0 1 14850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_184
timestamp 1675431861
transform 1 0 5500 0 1 15950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_185
timestamp 1675431861
transform 1 0 5500 0 1 17050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_186
timestamp 1675431861
transform 1 0 5500 0 1 18150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_187
timestamp 1675431861
transform 1 0 6050 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_188
timestamp 1675431861
transform 1 0 6050 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_189
timestamp 1675431861
transform 1 0 6050 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_190
timestamp 1675431861
transform 1 0 6050 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_191
timestamp 1675431861
transform 1 0 6050 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_192
timestamp 1675431861
transform 1 0 6050 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_193
timestamp 1675431861
transform 1 0 6050 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_194
timestamp 1675431861
transform 1 0 6050 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_195
timestamp 1675431861
transform 1 0 6050 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_196
timestamp 1675431861
transform 1 0 6050 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_197
timestamp 1675431861
transform 1 0 6050 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_198
timestamp 1675431861
transform 1 0 6050 0 1 12100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_199
timestamp 1675431861
transform 1 0 6050 0 1 13200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_200
timestamp 1675431861
transform 1 0 6050 0 1 14300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_201
timestamp 1675431861
transform 1 0 6050 0 1 15400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_202
timestamp 1675431861
transform 1 0 6050 0 1 16500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_203
timestamp 1675431861
transform 1 0 6050 0 1 17600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_204
timestamp 1675431861
transform 1 0 6600 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_205
timestamp 1675431861
transform 1 0 6600 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_206
timestamp 1675431861
transform 1 0 6600 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_207
timestamp 1675431861
transform 1 0 6600 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_208
timestamp 1675431861
transform 1 0 6600 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_209
timestamp 1675431861
transform 1 0 6600 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_210
timestamp 1675431861
transform 1 0 6600 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_211
timestamp 1675431861
transform 1 0 6600 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_212
timestamp 1675431861
transform 1 0 6600 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_213
timestamp 1675431861
transform 1 0 6600 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_214
timestamp 1675431861
transform 1 0 6600 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_215
timestamp 1675431861
transform 1 0 6600 0 1 12650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_216
timestamp 1675431861
transform 1 0 6600 0 1 13750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_217
timestamp 1675431861
transform 1 0 6600 0 1 14850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_218
timestamp 1675431861
transform 1 0 6600 0 1 15950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_219
timestamp 1675431861
transform 1 0 6600 0 1 17050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_220
timestamp 1675431861
transform 1 0 6600 0 1 18150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_221
timestamp 1675431861
transform 1 0 7150 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_222
timestamp 1675431861
transform 1 0 7150 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_223
timestamp 1675431861
transform 1 0 7150 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_224
timestamp 1675431861
transform 1 0 7150 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_225
timestamp 1675431861
transform 1 0 7150 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_226
timestamp 1675431861
transform 1 0 7150 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_227
timestamp 1675431861
transform 1 0 7150 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_228
timestamp 1675431861
transform 1 0 7150 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_229
timestamp 1675431861
transform 1 0 7150 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_230
timestamp 1675431861
transform 1 0 7150 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_231
timestamp 1675431861
transform 1 0 7150 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_232
timestamp 1675431861
transform 1 0 7150 0 1 12100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_233
timestamp 1675431861
transform 1 0 7150 0 1 13200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_234
timestamp 1675431861
transform 1 0 7150 0 1 14300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_235
timestamp 1675431861
transform 1 0 7150 0 1 15400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_236
timestamp 1675431861
transform 1 0 7150 0 1 16500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_237
timestamp 1675431861
transform 1 0 7150 0 1 17600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_238
timestamp 1675431861
transform 1 0 7700 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_239
timestamp 1675431861
transform 1 0 7700 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_240
timestamp 1675431861
transform 1 0 7700 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_241
timestamp 1675431861
transform 1 0 7700 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_242
timestamp 1675431861
transform 1 0 7700 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_243
timestamp 1675431861
transform 1 0 7700 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_244
timestamp 1675431861
transform 1 0 7700 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_245
timestamp 1675431861
transform 1 0 7700 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_246
timestamp 1675431861
transform 1 0 7700 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_247
timestamp 1675431861
transform 1 0 7700 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_248
timestamp 1675431861
transform 1 0 7700 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_249
timestamp 1675431861
transform 1 0 7700 0 1 12650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_250
timestamp 1675431861
transform 1 0 7700 0 1 13750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_251
timestamp 1675431861
transform 1 0 7700 0 1 14850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_252
timestamp 1675431861
transform 1 0 7700 0 1 15950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_253
timestamp 1675431861
transform 1 0 7700 0 1 17050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_254
timestamp 1675431861
transform 1 0 7700 0 1 18150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_255
timestamp 1675431861
transform 1 0 8250 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_256
timestamp 1675431861
transform 1 0 8250 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_257
timestamp 1675431861
transform 1 0 8250 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_258
timestamp 1675431861
transform 1 0 8250 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_259
timestamp 1675431861
transform 1 0 8250 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_260
timestamp 1675431861
transform 1 0 8250 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_261
timestamp 1675431861
transform 1 0 8250 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_262
timestamp 1675431861
transform 1 0 8250 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_263
timestamp 1675431861
transform 1 0 8250 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_264
timestamp 1675431861
transform 1 0 8250 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_265
timestamp 1675431861
transform 1 0 8250 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_266
timestamp 1675431861
transform 1 0 8250 0 1 12100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_267
timestamp 1675431861
transform 1 0 8250 0 1 13200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_268
timestamp 1675431861
transform 1 0 8250 0 1 14300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_269
timestamp 1675431861
transform 1 0 8250 0 1 15400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_270
timestamp 1675431861
transform 1 0 8250 0 1 16500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_271
timestamp 1675431861
transform 1 0 8250 0 1 17600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_272
timestamp 1675431861
transform 1 0 8800 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_273
timestamp 1675431861
transform 1 0 8800 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_274
timestamp 1675431861
transform 1 0 8800 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_275
timestamp 1675431861
transform 1 0 8800 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_276
timestamp 1675431861
transform 1 0 8800 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_277
timestamp 1675431861
transform 1 0 8800 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_278
timestamp 1675431861
transform 1 0 8800 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_279
timestamp 1675431861
transform 1 0 8800 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_280
timestamp 1675431861
transform 1 0 8800 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_281
timestamp 1675431861
transform 1 0 8800 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_282
timestamp 1675431861
transform 1 0 8800 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_283
timestamp 1675431861
transform 1 0 8800 0 1 12650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_284
timestamp 1675431861
transform 1 0 8800 0 1 13750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_285
timestamp 1675431861
transform 1 0 8800 0 1 14850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_286
timestamp 1675431861
transform 1 0 8800 0 1 15950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_287
timestamp 1675431861
transform 1 0 8800 0 1 17050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_288
timestamp 1675431861
transform 1 0 8800 0 1 18150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_289
timestamp 1675431861
transform 1 0 9350 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_290
timestamp 1675431861
transform 1 0 9350 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_291
timestamp 1675431861
transform 1 0 9350 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_292
timestamp 1675431861
transform 1 0 9350 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_293
timestamp 1675431861
transform 1 0 9350 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_294
timestamp 1675431861
transform 1 0 9350 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_295
timestamp 1675431861
transform 1 0 9350 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_296
timestamp 1675431861
transform 1 0 9350 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_297
timestamp 1675431861
transform 1 0 9350 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_298
timestamp 1675431861
transform 1 0 9350 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_299
timestamp 1675431861
transform 1 0 9350 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_300
timestamp 1675431861
transform 1 0 9350 0 1 12100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_301
timestamp 1675431861
transform 1 0 9350 0 1 13200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_302
timestamp 1675431861
transform 1 0 9350 0 1 14300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_303
timestamp 1675431861
transform 1 0 9350 0 1 15400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_304
timestamp 1675431861
transform 1 0 9350 0 1 16500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_305
timestamp 1675431861
transform 1 0 9350 0 1 17600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_306
timestamp 1675431861
transform 1 0 9900 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_307
timestamp 1675431861
transform 1 0 9900 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_308
timestamp 1675431861
transform 1 0 9900 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_309
timestamp 1675431861
transform 1 0 9900 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_310
timestamp 1675431861
transform 1 0 9900 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_311
timestamp 1675431861
transform 1 0 9900 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_312
timestamp 1675431861
transform 1 0 9900 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_313
timestamp 1675431861
transform 1 0 9900 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_314
timestamp 1675431861
transform 1 0 9900 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_315
timestamp 1675431861
transform 1 0 9900 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_316
timestamp 1675431861
transform 1 0 9900 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_317
timestamp 1675431861
transform 1 0 9900 0 1 12650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_318
timestamp 1675431861
transform 1 0 9900 0 1 13750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_319
timestamp 1675431861
transform 1 0 9900 0 1 14850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_320
timestamp 1675431861
transform 1 0 9900 0 1 15950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_321
timestamp 1675431861
transform 1 0 9900 0 1 17050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_322
timestamp 1675431861
transform 1 0 9900 0 1 18150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_323
timestamp 1675431861
transform 1 0 10450 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_324
timestamp 1675431861
transform 1 0 10450 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_325
timestamp 1675431861
transform 1 0 10450 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_326
timestamp 1675431861
transform 1 0 10450 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_327
timestamp 1675431861
transform 1 0 10450 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_328
timestamp 1675431861
transform 1 0 10450 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_329
timestamp 1675431861
transform 1 0 10450 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_330
timestamp 1675431861
transform 1 0 10450 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_331
timestamp 1675431861
transform 1 0 10450 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_332
timestamp 1675431861
transform 1 0 10450 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_333
timestamp 1675431861
transform 1 0 10450 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_334
timestamp 1675431861
transform 1 0 10450 0 1 12100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_335
timestamp 1675431861
transform 1 0 10450 0 1 13200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_336
timestamp 1675431861
transform 1 0 10450 0 1 14300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_337
timestamp 1675431861
transform 1 0 10450 0 1 15400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_338
timestamp 1675431861
transform 1 0 10450 0 1 16500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_339
timestamp 1675431861
transform 1 0 10450 0 1 17600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_340
timestamp 1675431861
transform 1 0 11000 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_341
timestamp 1675431861
transform 1 0 11000 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_342
timestamp 1675431861
transform 1 0 11000 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_343
timestamp 1675431861
transform 1 0 11000 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_344
timestamp 1675431861
transform 1 0 11000 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_345
timestamp 1675431861
transform 1 0 11000 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_346
timestamp 1675431861
transform 1 0 11000 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_347
timestamp 1675431861
transform 1 0 11000 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_348
timestamp 1675431861
transform 1 0 11000 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_349
timestamp 1675431861
transform 1 0 11000 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_350
timestamp 1675431861
transform 1 0 11000 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_351
timestamp 1675431861
transform 1 0 11000 0 1 12650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_352
timestamp 1675431861
transform 1 0 11000 0 1 13750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_353
timestamp 1675431861
transform 1 0 11000 0 1 14850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_354
timestamp 1675431861
transform 1 0 11000 0 1 15950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_355
timestamp 1675431861
transform 1 0 11000 0 1 17050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_356
timestamp 1675431861
transform 1 0 11000 0 1 18150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_357
timestamp 1675431861
transform 1 0 11550 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_358
timestamp 1675431861
transform 1 0 11550 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_359
timestamp 1675431861
transform 1 0 11550 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_360
timestamp 1675431861
transform 1 0 11550 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_361
timestamp 1675431861
transform 1 0 11550 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_362
timestamp 1675431861
transform 1 0 11550 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_363
timestamp 1675431861
transform 1 0 11550 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_364
timestamp 1675431861
transform 1 0 11550 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_365
timestamp 1675431861
transform 1 0 11550 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_366
timestamp 1675431861
transform 1 0 11550 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_367
timestamp 1675431861
transform 1 0 11550 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_368
timestamp 1675431861
transform 1 0 11550 0 1 12100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_369
timestamp 1675431861
transform 1 0 11550 0 1 13200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_370
timestamp 1675431861
transform 1 0 11550 0 1 14300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_371
timestamp 1675431861
transform 1 0 11550 0 1 15400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_372
timestamp 1675431861
transform 1 0 11550 0 1 16500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_373
timestamp 1675431861
transform 1 0 11550 0 1 17600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_374
timestamp 1675431861
transform 1 0 12100 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_375
timestamp 1675431861
transform 1 0 12100 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_376
timestamp 1675431861
transform 1 0 12100 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_377
timestamp 1675431861
transform 1 0 12100 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_378
timestamp 1675431861
transform 1 0 12100 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_379
timestamp 1675431861
transform 1 0 12100 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_380
timestamp 1675431861
transform 1 0 12100 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_381
timestamp 1675431861
transform 1 0 12100 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_382
timestamp 1675431861
transform 1 0 12100 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_383
timestamp 1675431861
transform 1 0 12100 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_384
timestamp 1675431861
transform 1 0 12100 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_385
timestamp 1675431861
transform 1 0 12100 0 1 12650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_386
timestamp 1675431861
transform 1 0 12100 0 1 13750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_387
timestamp 1675431861
transform 1 0 12100 0 1 14850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_388
timestamp 1675431861
transform 1 0 12100 0 1 15950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_389
timestamp 1675431861
transform 1 0 12100 0 1 17050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_390
timestamp 1675431861
transform 1 0 12100 0 1 18150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_391
timestamp 1675431861
transform 1 0 12650 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_392
timestamp 1675431861
transform 1 0 12650 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_393
timestamp 1675431861
transform 1 0 12650 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_394
timestamp 1675431861
transform 1 0 12650 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_395
timestamp 1675431861
transform 1 0 12650 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_396
timestamp 1675431861
transform 1 0 12650 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_397
timestamp 1675431861
transform 1 0 12650 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_398
timestamp 1675431861
transform 1 0 12650 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_399
timestamp 1675431861
transform 1 0 12650 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_400
timestamp 1675431861
transform 1 0 12650 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_401
timestamp 1675431861
transform 1 0 12650 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_402
timestamp 1675431861
transform 1 0 12650 0 1 12100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_403
timestamp 1675431861
transform 1 0 12650 0 1 13200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_404
timestamp 1675431861
transform 1 0 12650 0 1 14300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_405
timestamp 1675431861
transform 1 0 12650 0 1 15400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_406
timestamp 1675431861
transform 1 0 12650 0 1 16500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_407
timestamp 1675431861
transform 1 0 12650 0 1 17600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_408
timestamp 1675431861
transform 1 0 13200 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_409
timestamp 1675431861
transform 1 0 13200 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_410
timestamp 1675431861
transform 1 0 13200 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_411
timestamp 1675431861
transform 1 0 13200 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_412
timestamp 1675431861
transform 1 0 13200 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_413
timestamp 1675431861
transform 1 0 13200 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_414
timestamp 1675431861
transform 1 0 13200 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_415
timestamp 1675431861
transform 1 0 13200 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_416
timestamp 1675431861
transform 1 0 13200 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_417
timestamp 1675431861
transform 1 0 13200 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_418
timestamp 1675431861
transform 1 0 13200 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_419
timestamp 1675431861
transform 1 0 13200 0 1 12650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_420
timestamp 1675431861
transform 1 0 13200 0 1 13750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_421
timestamp 1675431861
transform 1 0 13200 0 1 14850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_422
timestamp 1675431861
transform 1 0 13200 0 1 15950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_423
timestamp 1675431861
transform 1 0 13200 0 1 17050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_424
timestamp 1675431861
transform 1 0 13200 0 1 18150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_425
timestamp 1675431861
transform 1 0 13750 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_426
timestamp 1675431861
transform 1 0 13750 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_427
timestamp 1675431861
transform 1 0 13750 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_428
timestamp 1675431861
transform 1 0 13750 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_429
timestamp 1675431861
transform 1 0 13750 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_430
timestamp 1675431861
transform 1 0 13750 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_431
timestamp 1675431861
transform 1 0 13750 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_432
timestamp 1675431861
transform 1 0 13750 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_433
timestamp 1675431861
transform 1 0 13750 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_434
timestamp 1675431861
transform 1 0 13750 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_435
timestamp 1675431861
transform 1 0 13750 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_436
timestamp 1675431861
transform 1 0 13750 0 1 12100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_437
timestamp 1675431861
transform 1 0 13750 0 1 13200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_438
timestamp 1675431861
transform 1 0 13750 0 1 14300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_439
timestamp 1675431861
transform 1 0 13750 0 1 15400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_440
timestamp 1675431861
transform 1 0 13750 0 1 16500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_441
timestamp 1675431861
transform 1 0 13750 0 1 17600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_442
timestamp 1675431861
transform 1 0 14300 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_443
timestamp 1675431861
transform 1 0 14300 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_444
timestamp 1675431861
transform 1 0 14300 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_445
timestamp 1675431861
transform 1 0 14300 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_446
timestamp 1675431861
transform 1 0 14300 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_447
timestamp 1675431861
transform 1 0 14300 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_448
timestamp 1675431861
transform 1 0 14300 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_449
timestamp 1675431861
transform 1 0 14300 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_450
timestamp 1675431861
transform 1 0 14300 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_451
timestamp 1675431861
transform 1 0 14300 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_452
timestamp 1675431861
transform 1 0 14300 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_453
timestamp 1675431861
transform 1 0 14300 0 1 12650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_454
timestamp 1675431861
transform 1 0 14300 0 1 13750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_455
timestamp 1675431861
transform 1 0 14300 0 1 14850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_456
timestamp 1675431861
transform 1 0 14300 0 1 15950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_457
timestamp 1675431861
transform 1 0 14300 0 1 17050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_458
timestamp 1675431861
transform 1 0 14300 0 1 18150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_459
timestamp 1675431861
transform 1 0 14850 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_460
timestamp 1675431861
transform 1 0 14850 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_461
timestamp 1675431861
transform 1 0 14850 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_462
timestamp 1675431861
transform 1 0 14850 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_463
timestamp 1675431861
transform 1 0 14850 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_464
timestamp 1675431861
transform 1 0 14850 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_465
timestamp 1675431861
transform 1 0 14850 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_466
timestamp 1675431861
transform 1 0 14850 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_467
timestamp 1675431861
transform 1 0 14850 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_468
timestamp 1675431861
transform 1 0 14850 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_469
timestamp 1675431861
transform 1 0 14850 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_470
timestamp 1675431861
transform 1 0 14850 0 1 12100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_471
timestamp 1675431861
transform 1 0 14850 0 1 13200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_472
timestamp 1675431861
transform 1 0 14850 0 1 14300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_473
timestamp 1675431861
transform 1 0 14850 0 1 15400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_474
timestamp 1675431861
transform 1 0 14850 0 1 16500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_475
timestamp 1675431861
transform 1 0 14850 0 1 17600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_476
timestamp 1675431861
transform 1 0 15400 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_477
timestamp 1675431861
transform 1 0 15400 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_478
timestamp 1675431861
transform 1 0 15400 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_479
timestamp 1675431861
transform 1 0 15400 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_480
timestamp 1675431861
transform 1 0 15400 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_481
timestamp 1675431861
transform 1 0 15400 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_482
timestamp 1675431861
transform 1 0 15400 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_483
timestamp 1675431861
transform 1 0 15400 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_484
timestamp 1675431861
transform 1 0 15400 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_485
timestamp 1675431861
transform 1 0 15400 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_486
timestamp 1675431861
transform 1 0 15400 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_487
timestamp 1675431861
transform 1 0 15400 0 1 12650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_488
timestamp 1675431861
transform 1 0 15400 0 1 13750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_489
timestamp 1675431861
transform 1 0 15400 0 1 14850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_490
timestamp 1675431861
transform 1 0 15400 0 1 15950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_491
timestamp 1675431861
transform 1 0 15400 0 1 17050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_492
timestamp 1675431861
transform 1 0 15400 0 1 18150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_493
timestamp 1675431861
transform 1 0 15950 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_494
timestamp 1675431861
transform 1 0 15950 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_495
timestamp 1675431861
transform 1 0 15950 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_496
timestamp 1675431861
transform 1 0 15950 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_497
timestamp 1675431861
transform 1 0 15950 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_498
timestamp 1675431861
transform 1 0 15950 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_499
timestamp 1675431861
transform 1 0 15950 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_500
timestamp 1675431861
transform 1 0 15950 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_501
timestamp 1675431861
transform 1 0 15950 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_502
timestamp 1675431861
transform 1 0 15950 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_503
timestamp 1675431861
transform 1 0 15950 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_504
timestamp 1675431861
transform 1 0 15950 0 1 12100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_505
timestamp 1675431861
transform 1 0 15950 0 1 13200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_506
timestamp 1675431861
transform 1 0 15950 0 1 14300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_507
timestamp 1675431861
transform 1 0 15950 0 1 15400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_508
timestamp 1675431861
transform 1 0 15950 0 1 16500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_509
timestamp 1675431861
transform 1 0 15950 0 1 17600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_510
timestamp 1675431861
transform 1 0 16500 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_511
timestamp 1675431861
transform 1 0 16500 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_512
timestamp 1675431861
transform 1 0 16500 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_513
timestamp 1675431861
transform 1 0 16500 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_514
timestamp 1675431861
transform 1 0 16500 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_515
timestamp 1675431861
transform 1 0 16500 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_516
timestamp 1675431861
transform 1 0 16500 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_517
timestamp 1675431861
transform 1 0 16500 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_518
timestamp 1675431861
transform 1 0 16500 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_519
timestamp 1675431861
transform 1 0 16500 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_520
timestamp 1675431861
transform 1 0 16500 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_521
timestamp 1675431861
transform 1 0 16500 0 1 12650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_522
timestamp 1675431861
transform 1 0 16500 0 1 13750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_523
timestamp 1675431861
transform 1 0 16500 0 1 14850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_524
timestamp 1675431861
transform 1 0 16500 0 1 15950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_525
timestamp 1675431861
transform 1 0 16500 0 1 17050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_526
timestamp 1675431861
transform 1 0 16500 0 1 18150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_527
timestamp 1675431861
transform 1 0 17050 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_528
timestamp 1675431861
transform 1 0 17050 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_529
timestamp 1675431861
transform 1 0 17050 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_530
timestamp 1675431861
transform 1 0 17050 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_531
timestamp 1675431861
transform 1 0 17050 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_532
timestamp 1675431861
transform 1 0 17050 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_533
timestamp 1675431861
transform 1 0 17050 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_534
timestamp 1675431861
transform 1 0 17050 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_535
timestamp 1675431861
transform 1 0 17050 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_536
timestamp 1675431861
transform 1 0 17050 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_537
timestamp 1675431861
transform 1 0 17050 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_538
timestamp 1675431861
transform 1 0 17050 0 1 12100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_539
timestamp 1675431861
transform 1 0 17050 0 1 13200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_540
timestamp 1675431861
transform 1 0 17050 0 1 14300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_541
timestamp 1675431861
transform 1 0 17050 0 1 15400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_542
timestamp 1675431861
transform 1 0 17050 0 1 16500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_543
timestamp 1675431861
transform 1 0 17050 0 1 17600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_544
timestamp 1675431861
transform 1 0 17600 0 1 550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_545
timestamp 1675431861
transform 1 0 17600 0 1 1650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_546
timestamp 1675431861
transform 1 0 17600 0 1 2750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_547
timestamp 1675431861
transform 1 0 17600 0 1 3850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_548
timestamp 1675431861
transform 1 0 17600 0 1 4950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_549
timestamp 1675431861
transform 1 0 17600 0 1 6050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_550
timestamp 1675431861
transform 1 0 17600 0 1 7150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_551
timestamp 1675431861
transform 1 0 17600 0 1 8250
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_552
timestamp 1675431861
transform 1 0 17600 0 1 9350
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_553
timestamp 1675431861
transform 1 0 17600 0 1 10450
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_554
timestamp 1675431861
transform 1 0 17600 0 1 11550
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_555
timestamp 1675431861
transform 1 0 17600 0 1 12650
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_556
timestamp 1675431861
transform 1 0 17600 0 1 13750
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_557
timestamp 1675431861
transform 1 0 17600 0 1 14850
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_558
timestamp 1675431861
transform 1 0 17600 0 1 15950
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_559
timestamp 1675431861
transform 1 0 17600 0 1 17050
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_560
timestamp 1675431861
transform 1 0 17600 0 1 18150
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_561
timestamp 1675431861
transform 1 0 18150 0 1 0
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_562
timestamp 1675431861
transform 1 0 18150 0 1 1100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_563
timestamp 1675431861
transform 1 0 18150 0 1 2200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_564
timestamp 1675431861
transform 1 0 18150 0 1 3300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_565
timestamp 1675431861
transform 1 0 18150 0 1 4400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_566
timestamp 1675431861
transform 1 0 18150 0 1 5500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_567
timestamp 1675431861
transform 1 0 18150 0 1 6600
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_568
timestamp 1675431861
transform 1 0 18150 0 1 7700
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_569
timestamp 1675431861
transform 1 0 18150 0 1 8800
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_570
timestamp 1675431861
transform 1 0 18150 0 1 9900
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_571
timestamp 1675431861
transform 1 0 18150 0 1 11000
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_572
timestamp 1675431861
transform 1 0 18150 0 1 12100
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_573
timestamp 1675431861
transform 1 0 18150 0 1 13200
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_574
timestamp 1675431861
transform 1 0 18150 0 1 14300
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_575
timestamp 1675431861
transform 1 0 18150 0 1 15400
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_576
timestamp 1675431861
transform 1 0 18150 0 1 16500
box -113 -113 663 663
use nmos_drain_in  nmos_drain_in_577
timestamp 1675431861
transform 1 0 18150 0 1 17600
box -113 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_0 waffle_cells
timestamp 1675431308
transform 0 -1 550 -1 0 19250
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_1
timestamp 1675431308
transform 1 0 -550 0 1 550
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_2
timestamp 1675431308
transform 0 -1 1650 -1 0 19250
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_3
timestamp 1675431308
transform 1 0 -550 0 1 1650
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_4
timestamp 1675431308
transform 0 -1 2750 -1 0 19250
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_5
timestamp 1675431308
transform 1 0 -550 0 1 2750
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_6
timestamp 1675431308
transform 0 -1 3850 -1 0 19250
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_7
timestamp 1675431308
transform 1 0 -550 0 1 3850
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_8
timestamp 1675431308
transform 0 -1 4950 -1 0 19250
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_9
timestamp 1675431308
transform 1 0 -550 0 1 4950
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_10
timestamp 1675431308
transform 0 -1 6050 -1 0 19250
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_11
timestamp 1675431308
transform 1 0 -550 0 1 6050
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_12
timestamp 1675431308
transform 0 -1 7150 -1 0 19250
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_13
timestamp 1675431308
transform 1 0 -550 0 1 7150
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_14
timestamp 1675431308
transform 0 -1 8250 -1 0 19250
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_15
timestamp 1675431308
transform 1 0 -550 0 1 8250
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_16
timestamp 1675431308
transform 0 -1 9350 -1 0 19250
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_17
timestamp 1675431308
transform 1 0 -550 0 1 9350
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_18
timestamp 1675431308
transform 0 -1 10450 -1 0 19250
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_19
timestamp 1675431308
transform 1 0 -550 0 1 10450
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_20
timestamp 1675431308
transform 0 -1 11550 -1 0 19250
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_21
timestamp 1675431308
transform 1 0 -550 0 1 11550
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_22
timestamp 1675431308
transform 0 -1 12650 -1 0 19250
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_23
timestamp 1675431308
transform 1 0 -550 0 1 12650
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_24
timestamp 1675431308
transform 0 -1 13750 -1 0 19250
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_25
timestamp 1675431308
transform 1 0 -550 0 1 13750
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_26
timestamp 1675431308
transform 0 -1 14850 -1 0 19250
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_27
timestamp 1675431308
transform 1 0 -550 0 1 14850
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_28
timestamp 1675431308
transform 0 -1 15950 -1 0 19250
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_29
timestamp 1675431308
transform 1 0 -550 0 1 15950
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_30
timestamp 1675431308
transform 0 -1 17050 -1 0 19250
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_31
timestamp 1675431308
transform 1 0 -550 0 1 17050
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_32
timestamp 1675431308
transform 0 -1 18150 -1 0 19250
box -975 -113 663 663
use nmos_source_frame_lt  nmos_source_frame_lt_33
timestamp 1675431308
transform 1 0 -550 0 1 18150
box -975 -113 663 663
use nmos_source_frame_rb  nmos_source_frame_rb_0 waffle_cells
timestamp 1675430904
transform 1 0 18700 0 1 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_1
timestamp 1675430904
transform 0 -1 1100 -1 0 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_2
timestamp 1675430904
transform 1 0 18700 0 1 1100
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_3
timestamp 1675430904
transform 0 -1 2200 -1 0 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_4
timestamp 1675430904
transform 1 0 18700 0 1 2200
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_5
timestamp 1675430904
transform 0 -1 3300 -1 0 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_6
timestamp 1675430904
transform 1 0 18700 0 1 3300
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_7
timestamp 1675430904
transform 0 -1 4400 -1 0 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_8
timestamp 1675430904
transform 1 0 18700 0 1 4400
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_9
timestamp 1675430904
transform 0 -1 5500 -1 0 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_10
timestamp 1675430904
transform 1 0 18700 0 1 5500
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_11
timestamp 1675430904
transform 0 -1 6600 -1 0 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_12
timestamp 1675430904
transform 1 0 18700 0 1 6600
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_13
timestamp 1675430904
transform 0 -1 7700 -1 0 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_14
timestamp 1675430904
transform 1 0 18700 0 1 7700
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_15
timestamp 1675430904
transform 0 -1 8800 -1 0 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_16
timestamp 1675430904
transform 1 0 18700 0 1 8800
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_17
timestamp 1675430904
transform 0 -1 9900 -1 0 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_18
timestamp 1675430904
transform 1 0 18700 0 1 9900
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_19
timestamp 1675430904
transform 0 -1 11000 -1 0 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_20
timestamp 1675430904
transform 1 0 18700 0 1 11000
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_21
timestamp 1675430904
transform 0 -1 12100 -1 0 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_22
timestamp 1675430904
transform 1 0 18700 0 1 12100
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_23
timestamp 1675430904
transform 0 -1 13200 -1 0 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_24
timestamp 1675430904
transform 1 0 18700 0 1 13200
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_25
timestamp 1675430904
transform 0 -1 14300 -1 0 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_26
timestamp 1675430904
transform 1 0 18700 0 1 14300
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_27
timestamp 1675430904
transform 0 -1 15400 -1 0 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_28
timestamp 1675430904
transform 1 0 18700 0 1 15400
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_29
timestamp 1675430904
transform 0 -1 16500 -1 0 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_30
timestamp 1675430904
transform 1 0 18700 0 1 16500
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_31
timestamp 1675430904
transform 0 -1 17600 -1 0 0
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_32
timestamp 1675430904
transform 1 0 18700 0 1 17600
box -113 -113 1575 663
use nmos_source_frame_rb  nmos_source_frame_rb_33
timestamp 1675430904
transform 0 -1 18700 -1 0 0
box -113 -113 1575 663
use nmos_source_in  nmos_source_in_0 waffle_cells
timestamp 1675431769
transform 1 0 0 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_1
timestamp 1675431769
transform 1 0 0 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_2
timestamp 1675431769
transform 1 0 0 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_3
timestamp 1675431769
transform 1 0 0 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_4
timestamp 1675431769
transform 1 0 0 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_5
timestamp 1675431769
transform 1 0 0 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_6
timestamp 1675431769
transform 1 0 0 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_7
timestamp 1675431769
transform 1 0 0 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_8
timestamp 1675431769
transform 1 0 0 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_9
timestamp 1675431769
transform 1 0 0 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_10
timestamp 1675431769
transform 1 0 0 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_11
timestamp 1675431769
transform 1 0 0 0 1 12100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_12
timestamp 1675431769
transform 1 0 0 0 1 13200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_13
timestamp 1675431769
transform 1 0 0 0 1 14300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_14
timestamp 1675431769
transform 1 0 0 0 1 15400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_15
timestamp 1675431769
transform 1 0 0 0 1 16500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_16
timestamp 1675431769
transform 1 0 0 0 1 17600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_17
timestamp 1675431769
transform 1 0 550 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_18
timestamp 1675431769
transform 1 0 550 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_19
timestamp 1675431769
transform 1 0 550 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_20
timestamp 1675431769
transform 1 0 550 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_21
timestamp 1675431769
transform 1 0 550 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_22
timestamp 1675431769
transform 1 0 550 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_23
timestamp 1675431769
transform 1 0 550 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_24
timestamp 1675431769
transform 1 0 550 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_25
timestamp 1675431769
transform 1 0 550 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_26
timestamp 1675431769
transform 1 0 550 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_27
timestamp 1675431769
transform 1 0 550 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_28
timestamp 1675431769
transform 1 0 550 0 1 12650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_29
timestamp 1675431769
transform 1 0 550 0 1 13750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_30
timestamp 1675431769
transform 1 0 550 0 1 14850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_31
timestamp 1675431769
transform 1 0 550 0 1 15950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_32
timestamp 1675431769
transform 1 0 550 0 1 17050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_33
timestamp 1675431769
transform 1 0 550 0 1 18150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_34
timestamp 1675431769
transform 1 0 1100 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_35
timestamp 1675431769
transform 1 0 1100 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_36
timestamp 1675431769
transform 1 0 1100 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_37
timestamp 1675431769
transform 1 0 1100 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_38
timestamp 1675431769
transform 1 0 1100 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_39
timestamp 1675431769
transform 1 0 1100 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_40
timestamp 1675431769
transform 1 0 1100 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_41
timestamp 1675431769
transform 1 0 1100 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_42
timestamp 1675431769
transform 1 0 1100 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_43
timestamp 1675431769
transform 1 0 1100 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_44
timestamp 1675431769
transform 1 0 1100 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_45
timestamp 1675431769
transform 1 0 1100 0 1 12100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_46
timestamp 1675431769
transform 1 0 1100 0 1 13200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_47
timestamp 1675431769
transform 1 0 1100 0 1 14300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_48
timestamp 1675431769
transform 1 0 1100 0 1 15400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_49
timestamp 1675431769
transform 1 0 1100 0 1 16500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_50
timestamp 1675431769
transform 1 0 1100 0 1 17600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_51
timestamp 1675431769
transform 1 0 1650 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_52
timestamp 1675431769
transform 1 0 1650 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_53
timestamp 1675431769
transform 1 0 1650 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_54
timestamp 1675431769
transform 1 0 1650 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_55
timestamp 1675431769
transform 1 0 1650 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_56
timestamp 1675431769
transform 1 0 1650 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_57
timestamp 1675431769
transform 1 0 1650 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_58
timestamp 1675431769
transform 1 0 1650 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_59
timestamp 1675431769
transform 1 0 1650 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_60
timestamp 1675431769
transform 1 0 1650 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_61
timestamp 1675431769
transform 1 0 1650 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_62
timestamp 1675431769
transform 1 0 1650 0 1 12650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_63
timestamp 1675431769
transform 1 0 1650 0 1 13750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_64
timestamp 1675431769
transform 1 0 1650 0 1 14850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_65
timestamp 1675431769
transform 1 0 1650 0 1 15950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_66
timestamp 1675431769
transform 1 0 1650 0 1 17050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_67
timestamp 1675431769
transform 1 0 1650 0 1 18150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_68
timestamp 1675431769
transform 1 0 2200 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_69
timestamp 1675431769
transform 1 0 2200 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_70
timestamp 1675431769
transform 1 0 2200 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_71
timestamp 1675431769
transform 1 0 2200 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_72
timestamp 1675431769
transform 1 0 2200 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_73
timestamp 1675431769
transform 1 0 2200 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_74
timestamp 1675431769
transform 1 0 2200 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_75
timestamp 1675431769
transform 1 0 2200 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_76
timestamp 1675431769
transform 1 0 2200 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_77
timestamp 1675431769
transform 1 0 2200 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_78
timestamp 1675431769
transform 1 0 2200 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_79
timestamp 1675431769
transform 1 0 2200 0 1 12100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_80
timestamp 1675431769
transform 1 0 2200 0 1 13200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_81
timestamp 1675431769
transform 1 0 2200 0 1 14300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_82
timestamp 1675431769
transform 1 0 2200 0 1 15400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_83
timestamp 1675431769
transform 1 0 2200 0 1 16500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_84
timestamp 1675431769
transform 1 0 2200 0 1 17600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_85
timestamp 1675431769
transform 1 0 2750 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_86
timestamp 1675431769
transform 1 0 2750 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_87
timestamp 1675431769
transform 1 0 2750 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_88
timestamp 1675431769
transform 1 0 2750 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_89
timestamp 1675431769
transform 1 0 2750 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_90
timestamp 1675431769
transform 1 0 2750 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_91
timestamp 1675431769
transform 1 0 2750 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_92
timestamp 1675431769
transform 1 0 2750 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_93
timestamp 1675431769
transform 1 0 2750 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_94
timestamp 1675431769
transform 1 0 2750 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_95
timestamp 1675431769
transform 1 0 2750 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_96
timestamp 1675431769
transform 1 0 2750 0 1 12650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_97
timestamp 1675431769
transform 1 0 2750 0 1 13750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_98
timestamp 1675431769
transform 1 0 2750 0 1 14850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_99
timestamp 1675431769
transform 1 0 2750 0 1 15950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_100
timestamp 1675431769
transform 1 0 2750 0 1 17050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_101
timestamp 1675431769
transform 1 0 2750 0 1 18150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_102
timestamp 1675431769
transform 1 0 3300 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_103
timestamp 1675431769
transform 1 0 3300 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_104
timestamp 1675431769
transform 1 0 3300 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_105
timestamp 1675431769
transform 1 0 3300 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_106
timestamp 1675431769
transform 1 0 3300 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_107
timestamp 1675431769
transform 1 0 3300 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_108
timestamp 1675431769
transform 1 0 3300 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_109
timestamp 1675431769
transform 1 0 3300 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_110
timestamp 1675431769
transform 1 0 3300 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_111
timestamp 1675431769
transform 1 0 3300 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_112
timestamp 1675431769
transform 1 0 3300 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_113
timestamp 1675431769
transform 1 0 3300 0 1 12100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_114
timestamp 1675431769
transform 1 0 3300 0 1 13200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_115
timestamp 1675431769
transform 1 0 3300 0 1 14300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_116
timestamp 1675431769
transform 1 0 3300 0 1 15400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_117
timestamp 1675431769
transform 1 0 3300 0 1 16500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_118
timestamp 1675431769
transform 1 0 3300 0 1 17600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_119
timestamp 1675431769
transform 1 0 3850 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_120
timestamp 1675431769
transform 1 0 3850 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_121
timestamp 1675431769
transform 1 0 3850 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_122
timestamp 1675431769
transform 1 0 3850 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_123
timestamp 1675431769
transform 1 0 3850 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_124
timestamp 1675431769
transform 1 0 3850 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_125
timestamp 1675431769
transform 1 0 3850 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_126
timestamp 1675431769
transform 1 0 3850 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_127
timestamp 1675431769
transform 1 0 3850 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_128
timestamp 1675431769
transform 1 0 3850 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_129
timestamp 1675431769
transform 1 0 3850 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_130
timestamp 1675431769
transform 1 0 3850 0 1 12650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_131
timestamp 1675431769
transform 1 0 3850 0 1 13750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_132
timestamp 1675431769
transform 1 0 3850 0 1 14850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_133
timestamp 1675431769
transform 1 0 3850 0 1 15950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_134
timestamp 1675431769
transform 1 0 3850 0 1 17050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_135
timestamp 1675431769
transform 1 0 3850 0 1 18150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_136
timestamp 1675431769
transform 1 0 4400 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_137
timestamp 1675431769
transform 1 0 4400 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_138
timestamp 1675431769
transform 1 0 4400 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_139
timestamp 1675431769
transform 1 0 4400 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_140
timestamp 1675431769
transform 1 0 4400 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_141
timestamp 1675431769
transform 1 0 4400 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_142
timestamp 1675431769
transform 1 0 4400 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_143
timestamp 1675431769
transform 1 0 4400 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_144
timestamp 1675431769
transform 1 0 4400 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_145
timestamp 1675431769
transform 1 0 4400 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_146
timestamp 1675431769
transform 1 0 4400 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_147
timestamp 1675431769
transform 1 0 4400 0 1 12100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_148
timestamp 1675431769
transform 1 0 4400 0 1 13200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_149
timestamp 1675431769
transform 1 0 4400 0 1 14300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_150
timestamp 1675431769
transform 1 0 4400 0 1 15400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_151
timestamp 1675431769
transform 1 0 4400 0 1 16500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_152
timestamp 1675431769
transform 1 0 4400 0 1 17600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_153
timestamp 1675431769
transform 1 0 4950 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_154
timestamp 1675431769
transform 1 0 4950 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_155
timestamp 1675431769
transform 1 0 4950 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_156
timestamp 1675431769
transform 1 0 4950 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_157
timestamp 1675431769
transform 1 0 4950 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_158
timestamp 1675431769
transform 1 0 4950 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_159
timestamp 1675431769
transform 1 0 4950 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_160
timestamp 1675431769
transform 1 0 4950 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_161
timestamp 1675431769
transform 1 0 4950 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_162
timestamp 1675431769
transform 1 0 4950 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_163
timestamp 1675431769
transform 1 0 4950 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_164
timestamp 1675431769
transform 1 0 4950 0 1 12650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_165
timestamp 1675431769
transform 1 0 4950 0 1 13750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_166
timestamp 1675431769
transform 1 0 4950 0 1 14850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_167
timestamp 1675431769
transform 1 0 4950 0 1 15950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_168
timestamp 1675431769
transform 1 0 4950 0 1 17050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_169
timestamp 1675431769
transform 1 0 4950 0 1 18150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_170
timestamp 1675431769
transform 1 0 5500 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_171
timestamp 1675431769
transform 1 0 5500 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_172
timestamp 1675431769
transform 1 0 5500 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_173
timestamp 1675431769
transform 1 0 5500 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_174
timestamp 1675431769
transform 1 0 5500 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_175
timestamp 1675431769
transform 1 0 5500 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_176
timestamp 1675431769
transform 1 0 5500 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_177
timestamp 1675431769
transform 1 0 5500 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_178
timestamp 1675431769
transform 1 0 5500 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_179
timestamp 1675431769
transform 1 0 5500 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_180
timestamp 1675431769
transform 1 0 5500 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_181
timestamp 1675431769
transform 1 0 5500 0 1 12100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_182
timestamp 1675431769
transform 1 0 5500 0 1 13200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_183
timestamp 1675431769
transform 1 0 5500 0 1 14300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_184
timestamp 1675431769
transform 1 0 5500 0 1 15400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_185
timestamp 1675431769
transform 1 0 5500 0 1 16500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_186
timestamp 1675431769
transform 1 0 5500 0 1 17600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_187
timestamp 1675431769
transform 1 0 6050 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_188
timestamp 1675431769
transform 1 0 6050 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_189
timestamp 1675431769
transform 1 0 6050 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_190
timestamp 1675431769
transform 1 0 6050 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_191
timestamp 1675431769
transform 1 0 6050 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_192
timestamp 1675431769
transform 1 0 6050 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_193
timestamp 1675431769
transform 1 0 6050 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_194
timestamp 1675431769
transform 1 0 6050 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_195
timestamp 1675431769
transform 1 0 6050 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_196
timestamp 1675431769
transform 1 0 6050 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_197
timestamp 1675431769
transform 1 0 6050 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_198
timestamp 1675431769
transform 1 0 6050 0 1 12650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_199
timestamp 1675431769
transform 1 0 6050 0 1 13750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_200
timestamp 1675431769
transform 1 0 6050 0 1 14850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_201
timestamp 1675431769
transform 1 0 6050 0 1 15950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_202
timestamp 1675431769
transform 1 0 6050 0 1 17050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_203
timestamp 1675431769
transform 1 0 6050 0 1 18150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_204
timestamp 1675431769
transform 1 0 6600 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_205
timestamp 1675431769
transform 1 0 6600 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_206
timestamp 1675431769
transform 1 0 6600 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_207
timestamp 1675431769
transform 1 0 6600 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_208
timestamp 1675431769
transform 1 0 6600 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_209
timestamp 1675431769
transform 1 0 6600 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_210
timestamp 1675431769
transform 1 0 6600 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_211
timestamp 1675431769
transform 1 0 6600 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_212
timestamp 1675431769
transform 1 0 6600 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_213
timestamp 1675431769
transform 1 0 6600 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_214
timestamp 1675431769
transform 1 0 6600 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_215
timestamp 1675431769
transform 1 0 6600 0 1 12100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_216
timestamp 1675431769
transform 1 0 6600 0 1 13200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_217
timestamp 1675431769
transform 1 0 6600 0 1 14300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_218
timestamp 1675431769
transform 1 0 6600 0 1 15400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_219
timestamp 1675431769
transform 1 0 6600 0 1 16500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_220
timestamp 1675431769
transform 1 0 6600 0 1 17600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_221
timestamp 1675431769
transform 1 0 7150 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_222
timestamp 1675431769
transform 1 0 7150 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_223
timestamp 1675431769
transform 1 0 7150 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_224
timestamp 1675431769
transform 1 0 7150 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_225
timestamp 1675431769
transform 1 0 7150 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_226
timestamp 1675431769
transform 1 0 7150 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_227
timestamp 1675431769
transform 1 0 7150 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_228
timestamp 1675431769
transform 1 0 7150 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_229
timestamp 1675431769
transform 1 0 7150 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_230
timestamp 1675431769
transform 1 0 7150 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_231
timestamp 1675431769
transform 1 0 7150 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_232
timestamp 1675431769
transform 1 0 7150 0 1 12650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_233
timestamp 1675431769
transform 1 0 7150 0 1 13750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_234
timestamp 1675431769
transform 1 0 7150 0 1 14850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_235
timestamp 1675431769
transform 1 0 7150 0 1 15950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_236
timestamp 1675431769
transform 1 0 7150 0 1 17050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_237
timestamp 1675431769
transform 1 0 7150 0 1 18150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_238
timestamp 1675431769
transform 1 0 7700 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_239
timestamp 1675431769
transform 1 0 7700 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_240
timestamp 1675431769
transform 1 0 7700 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_241
timestamp 1675431769
transform 1 0 7700 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_242
timestamp 1675431769
transform 1 0 7700 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_243
timestamp 1675431769
transform 1 0 7700 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_244
timestamp 1675431769
transform 1 0 7700 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_245
timestamp 1675431769
transform 1 0 7700 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_246
timestamp 1675431769
transform 1 0 7700 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_247
timestamp 1675431769
transform 1 0 7700 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_248
timestamp 1675431769
transform 1 0 7700 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_249
timestamp 1675431769
transform 1 0 7700 0 1 12100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_250
timestamp 1675431769
transform 1 0 7700 0 1 13200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_251
timestamp 1675431769
transform 1 0 7700 0 1 14300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_252
timestamp 1675431769
transform 1 0 7700 0 1 15400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_253
timestamp 1675431769
transform 1 0 7700 0 1 16500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_254
timestamp 1675431769
transform 1 0 7700 0 1 17600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_255
timestamp 1675431769
transform 1 0 8250 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_256
timestamp 1675431769
transform 1 0 8250 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_257
timestamp 1675431769
transform 1 0 8250 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_258
timestamp 1675431769
transform 1 0 8250 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_259
timestamp 1675431769
transform 1 0 8250 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_260
timestamp 1675431769
transform 1 0 8250 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_261
timestamp 1675431769
transform 1 0 8250 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_262
timestamp 1675431769
transform 1 0 8250 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_263
timestamp 1675431769
transform 1 0 8250 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_264
timestamp 1675431769
transform 1 0 8250 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_265
timestamp 1675431769
transform 1 0 8250 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_266
timestamp 1675431769
transform 1 0 8250 0 1 12650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_267
timestamp 1675431769
transform 1 0 8250 0 1 13750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_268
timestamp 1675431769
transform 1 0 8250 0 1 14850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_269
timestamp 1675431769
transform 1 0 8250 0 1 15950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_270
timestamp 1675431769
transform 1 0 8250 0 1 17050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_271
timestamp 1675431769
transform 1 0 8250 0 1 18150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_272
timestamp 1675431769
transform 1 0 8800 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_273
timestamp 1675431769
transform 1 0 8800 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_274
timestamp 1675431769
transform 1 0 8800 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_275
timestamp 1675431769
transform 1 0 8800 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_276
timestamp 1675431769
transform 1 0 8800 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_277
timestamp 1675431769
transform 1 0 8800 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_278
timestamp 1675431769
transform 1 0 8800 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_279
timestamp 1675431769
transform 1 0 8800 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_280
timestamp 1675431769
transform 1 0 8800 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_281
timestamp 1675431769
transform 1 0 8800 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_282
timestamp 1675431769
transform 1 0 8800 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_283
timestamp 1675431769
transform 1 0 8800 0 1 12100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_284
timestamp 1675431769
transform 1 0 8800 0 1 13200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_285
timestamp 1675431769
transform 1 0 8800 0 1 14300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_286
timestamp 1675431769
transform 1 0 8800 0 1 15400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_287
timestamp 1675431769
transform 1 0 8800 0 1 16500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_288
timestamp 1675431769
transform 1 0 8800 0 1 17600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_289
timestamp 1675431769
transform 1 0 9350 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_290
timestamp 1675431769
transform 1 0 9350 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_291
timestamp 1675431769
transform 1 0 9350 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_292
timestamp 1675431769
transform 1 0 9350 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_293
timestamp 1675431769
transform 1 0 9350 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_294
timestamp 1675431769
transform 1 0 9350 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_295
timestamp 1675431769
transform 1 0 9350 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_296
timestamp 1675431769
transform 1 0 9350 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_297
timestamp 1675431769
transform 1 0 9350 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_298
timestamp 1675431769
transform 1 0 9350 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_299
timestamp 1675431769
transform 1 0 9350 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_300
timestamp 1675431769
transform 1 0 9350 0 1 12650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_301
timestamp 1675431769
transform 1 0 9350 0 1 13750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_302
timestamp 1675431769
transform 1 0 9350 0 1 14850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_303
timestamp 1675431769
transform 1 0 9350 0 1 15950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_304
timestamp 1675431769
transform 1 0 9350 0 1 17050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_305
timestamp 1675431769
transform 1 0 9350 0 1 18150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_306
timestamp 1675431769
transform 1 0 9900 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_307
timestamp 1675431769
transform 1 0 9900 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_308
timestamp 1675431769
transform 1 0 9900 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_309
timestamp 1675431769
transform 1 0 9900 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_310
timestamp 1675431769
transform 1 0 9900 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_311
timestamp 1675431769
transform 1 0 9900 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_312
timestamp 1675431769
transform 1 0 9900 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_313
timestamp 1675431769
transform 1 0 9900 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_314
timestamp 1675431769
transform 1 0 9900 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_315
timestamp 1675431769
transform 1 0 9900 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_316
timestamp 1675431769
transform 1 0 9900 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_317
timestamp 1675431769
transform 1 0 9900 0 1 12100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_318
timestamp 1675431769
transform 1 0 9900 0 1 13200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_319
timestamp 1675431769
transform 1 0 9900 0 1 14300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_320
timestamp 1675431769
transform 1 0 9900 0 1 15400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_321
timestamp 1675431769
transform 1 0 9900 0 1 16500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_322
timestamp 1675431769
transform 1 0 9900 0 1 17600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_323
timestamp 1675431769
transform 1 0 10450 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_324
timestamp 1675431769
transform 1 0 10450 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_325
timestamp 1675431769
transform 1 0 10450 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_326
timestamp 1675431769
transform 1 0 10450 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_327
timestamp 1675431769
transform 1 0 10450 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_328
timestamp 1675431769
transform 1 0 10450 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_329
timestamp 1675431769
transform 1 0 10450 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_330
timestamp 1675431769
transform 1 0 10450 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_331
timestamp 1675431769
transform 1 0 10450 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_332
timestamp 1675431769
transform 1 0 10450 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_333
timestamp 1675431769
transform 1 0 10450 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_334
timestamp 1675431769
transform 1 0 10450 0 1 12650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_335
timestamp 1675431769
transform 1 0 10450 0 1 13750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_336
timestamp 1675431769
transform 1 0 10450 0 1 14850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_337
timestamp 1675431769
transform 1 0 10450 0 1 15950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_338
timestamp 1675431769
transform 1 0 10450 0 1 17050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_339
timestamp 1675431769
transform 1 0 10450 0 1 18150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_340
timestamp 1675431769
transform 1 0 11000 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_341
timestamp 1675431769
transform 1 0 11000 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_342
timestamp 1675431769
transform 1 0 11000 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_343
timestamp 1675431769
transform 1 0 11000 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_344
timestamp 1675431769
transform 1 0 11000 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_345
timestamp 1675431769
transform 1 0 11000 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_346
timestamp 1675431769
transform 1 0 11000 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_347
timestamp 1675431769
transform 1 0 11000 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_348
timestamp 1675431769
transform 1 0 11000 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_349
timestamp 1675431769
transform 1 0 11000 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_350
timestamp 1675431769
transform 1 0 11000 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_351
timestamp 1675431769
transform 1 0 11000 0 1 12100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_352
timestamp 1675431769
transform 1 0 11000 0 1 13200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_353
timestamp 1675431769
transform 1 0 11000 0 1 14300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_354
timestamp 1675431769
transform 1 0 11000 0 1 15400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_355
timestamp 1675431769
transform 1 0 11000 0 1 16500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_356
timestamp 1675431769
transform 1 0 11000 0 1 17600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_357
timestamp 1675431769
transform 1 0 11550 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_358
timestamp 1675431769
transform 1 0 11550 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_359
timestamp 1675431769
transform 1 0 11550 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_360
timestamp 1675431769
transform 1 0 11550 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_361
timestamp 1675431769
transform 1 0 11550 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_362
timestamp 1675431769
transform 1 0 11550 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_363
timestamp 1675431769
transform 1 0 11550 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_364
timestamp 1675431769
transform 1 0 11550 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_365
timestamp 1675431769
transform 1 0 11550 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_366
timestamp 1675431769
transform 1 0 11550 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_367
timestamp 1675431769
transform 1 0 11550 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_368
timestamp 1675431769
transform 1 0 11550 0 1 12650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_369
timestamp 1675431769
transform 1 0 11550 0 1 13750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_370
timestamp 1675431769
transform 1 0 11550 0 1 14850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_371
timestamp 1675431769
transform 1 0 11550 0 1 15950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_372
timestamp 1675431769
transform 1 0 11550 0 1 17050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_373
timestamp 1675431769
transform 1 0 11550 0 1 18150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_374
timestamp 1675431769
transform 1 0 12100 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_375
timestamp 1675431769
transform 1 0 12100 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_376
timestamp 1675431769
transform 1 0 12100 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_377
timestamp 1675431769
transform 1 0 12100 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_378
timestamp 1675431769
transform 1 0 12100 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_379
timestamp 1675431769
transform 1 0 12100 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_380
timestamp 1675431769
transform 1 0 12100 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_381
timestamp 1675431769
transform 1 0 12100 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_382
timestamp 1675431769
transform 1 0 12100 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_383
timestamp 1675431769
transform 1 0 12100 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_384
timestamp 1675431769
transform 1 0 12100 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_385
timestamp 1675431769
transform 1 0 12100 0 1 12100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_386
timestamp 1675431769
transform 1 0 12100 0 1 13200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_387
timestamp 1675431769
transform 1 0 12100 0 1 14300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_388
timestamp 1675431769
transform 1 0 12100 0 1 15400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_389
timestamp 1675431769
transform 1 0 12100 0 1 16500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_390
timestamp 1675431769
transform 1 0 12100 0 1 17600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_391
timestamp 1675431769
transform 1 0 12650 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_392
timestamp 1675431769
transform 1 0 12650 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_393
timestamp 1675431769
transform 1 0 12650 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_394
timestamp 1675431769
transform 1 0 12650 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_395
timestamp 1675431769
transform 1 0 12650 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_396
timestamp 1675431769
transform 1 0 12650 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_397
timestamp 1675431769
transform 1 0 12650 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_398
timestamp 1675431769
transform 1 0 12650 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_399
timestamp 1675431769
transform 1 0 12650 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_400
timestamp 1675431769
transform 1 0 12650 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_401
timestamp 1675431769
transform 1 0 12650 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_402
timestamp 1675431769
transform 1 0 12650 0 1 12650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_403
timestamp 1675431769
transform 1 0 12650 0 1 13750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_404
timestamp 1675431769
transform 1 0 12650 0 1 14850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_405
timestamp 1675431769
transform 1 0 12650 0 1 15950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_406
timestamp 1675431769
transform 1 0 12650 0 1 17050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_407
timestamp 1675431769
transform 1 0 12650 0 1 18150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_408
timestamp 1675431769
transform 1 0 13200 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_409
timestamp 1675431769
transform 1 0 13200 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_410
timestamp 1675431769
transform 1 0 13200 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_411
timestamp 1675431769
transform 1 0 13200 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_412
timestamp 1675431769
transform 1 0 13200 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_413
timestamp 1675431769
transform 1 0 13200 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_414
timestamp 1675431769
transform 1 0 13200 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_415
timestamp 1675431769
transform 1 0 13200 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_416
timestamp 1675431769
transform 1 0 13200 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_417
timestamp 1675431769
transform 1 0 13200 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_418
timestamp 1675431769
transform 1 0 13200 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_419
timestamp 1675431769
transform 1 0 13200 0 1 12100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_420
timestamp 1675431769
transform 1 0 13200 0 1 13200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_421
timestamp 1675431769
transform 1 0 13200 0 1 14300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_422
timestamp 1675431769
transform 1 0 13200 0 1 15400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_423
timestamp 1675431769
transform 1 0 13200 0 1 16500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_424
timestamp 1675431769
transform 1 0 13200 0 1 17600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_425
timestamp 1675431769
transform 1 0 13750 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_426
timestamp 1675431769
transform 1 0 13750 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_427
timestamp 1675431769
transform 1 0 13750 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_428
timestamp 1675431769
transform 1 0 13750 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_429
timestamp 1675431769
transform 1 0 13750 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_430
timestamp 1675431769
transform 1 0 13750 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_431
timestamp 1675431769
transform 1 0 13750 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_432
timestamp 1675431769
transform 1 0 13750 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_433
timestamp 1675431769
transform 1 0 13750 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_434
timestamp 1675431769
transform 1 0 13750 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_435
timestamp 1675431769
transform 1 0 13750 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_436
timestamp 1675431769
transform 1 0 13750 0 1 12650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_437
timestamp 1675431769
transform 1 0 13750 0 1 13750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_438
timestamp 1675431769
transform 1 0 13750 0 1 14850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_439
timestamp 1675431769
transform 1 0 13750 0 1 15950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_440
timestamp 1675431769
transform 1 0 13750 0 1 17050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_441
timestamp 1675431769
transform 1 0 13750 0 1 18150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_442
timestamp 1675431769
transform 1 0 14300 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_443
timestamp 1675431769
transform 1 0 14300 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_444
timestamp 1675431769
transform 1 0 14300 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_445
timestamp 1675431769
transform 1 0 14300 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_446
timestamp 1675431769
transform 1 0 14300 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_447
timestamp 1675431769
transform 1 0 14300 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_448
timestamp 1675431769
transform 1 0 14300 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_449
timestamp 1675431769
transform 1 0 14300 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_450
timestamp 1675431769
transform 1 0 14300 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_451
timestamp 1675431769
transform 1 0 14300 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_452
timestamp 1675431769
transform 1 0 14300 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_453
timestamp 1675431769
transform 1 0 14300 0 1 12100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_454
timestamp 1675431769
transform 1 0 14300 0 1 13200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_455
timestamp 1675431769
transform 1 0 14300 0 1 14300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_456
timestamp 1675431769
transform 1 0 14300 0 1 15400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_457
timestamp 1675431769
transform 1 0 14300 0 1 16500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_458
timestamp 1675431769
transform 1 0 14300 0 1 17600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_459
timestamp 1675431769
transform 1 0 14850 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_460
timestamp 1675431769
transform 1 0 14850 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_461
timestamp 1675431769
transform 1 0 14850 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_462
timestamp 1675431769
transform 1 0 14850 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_463
timestamp 1675431769
transform 1 0 14850 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_464
timestamp 1675431769
transform 1 0 14850 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_465
timestamp 1675431769
transform 1 0 14850 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_466
timestamp 1675431769
transform 1 0 14850 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_467
timestamp 1675431769
transform 1 0 14850 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_468
timestamp 1675431769
transform 1 0 14850 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_469
timestamp 1675431769
transform 1 0 14850 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_470
timestamp 1675431769
transform 1 0 14850 0 1 12650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_471
timestamp 1675431769
transform 1 0 14850 0 1 13750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_472
timestamp 1675431769
transform 1 0 14850 0 1 14850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_473
timestamp 1675431769
transform 1 0 14850 0 1 15950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_474
timestamp 1675431769
transform 1 0 14850 0 1 17050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_475
timestamp 1675431769
transform 1 0 14850 0 1 18150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_476
timestamp 1675431769
transform 1 0 15400 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_477
timestamp 1675431769
transform 1 0 15400 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_478
timestamp 1675431769
transform 1 0 15400 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_479
timestamp 1675431769
transform 1 0 15400 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_480
timestamp 1675431769
transform 1 0 15400 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_481
timestamp 1675431769
transform 1 0 15400 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_482
timestamp 1675431769
transform 1 0 15400 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_483
timestamp 1675431769
transform 1 0 15400 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_484
timestamp 1675431769
transform 1 0 15400 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_485
timestamp 1675431769
transform 1 0 15400 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_486
timestamp 1675431769
transform 1 0 15400 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_487
timestamp 1675431769
transform 1 0 15400 0 1 12100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_488
timestamp 1675431769
transform 1 0 15400 0 1 13200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_489
timestamp 1675431769
transform 1 0 15400 0 1 14300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_490
timestamp 1675431769
transform 1 0 15400 0 1 15400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_491
timestamp 1675431769
transform 1 0 15400 0 1 16500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_492
timestamp 1675431769
transform 1 0 15400 0 1 17600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_493
timestamp 1675431769
transform 1 0 15950 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_494
timestamp 1675431769
transform 1 0 15950 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_495
timestamp 1675431769
transform 1 0 15950 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_496
timestamp 1675431769
transform 1 0 15950 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_497
timestamp 1675431769
transform 1 0 15950 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_498
timestamp 1675431769
transform 1 0 15950 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_499
timestamp 1675431769
transform 1 0 15950 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_500
timestamp 1675431769
transform 1 0 15950 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_501
timestamp 1675431769
transform 1 0 15950 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_502
timestamp 1675431769
transform 1 0 15950 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_503
timestamp 1675431769
transform 1 0 15950 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_504
timestamp 1675431769
transform 1 0 15950 0 1 12650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_505
timestamp 1675431769
transform 1 0 15950 0 1 13750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_506
timestamp 1675431769
transform 1 0 15950 0 1 14850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_507
timestamp 1675431769
transform 1 0 15950 0 1 15950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_508
timestamp 1675431769
transform 1 0 15950 0 1 17050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_509
timestamp 1675431769
transform 1 0 15950 0 1 18150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_510
timestamp 1675431769
transform 1 0 16500 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_511
timestamp 1675431769
transform 1 0 16500 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_512
timestamp 1675431769
transform 1 0 16500 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_513
timestamp 1675431769
transform 1 0 16500 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_514
timestamp 1675431769
transform 1 0 16500 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_515
timestamp 1675431769
transform 1 0 16500 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_516
timestamp 1675431769
transform 1 0 16500 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_517
timestamp 1675431769
transform 1 0 16500 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_518
timestamp 1675431769
transform 1 0 16500 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_519
timestamp 1675431769
transform 1 0 16500 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_520
timestamp 1675431769
transform 1 0 16500 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_521
timestamp 1675431769
transform 1 0 16500 0 1 12100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_522
timestamp 1675431769
transform 1 0 16500 0 1 13200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_523
timestamp 1675431769
transform 1 0 16500 0 1 14300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_524
timestamp 1675431769
transform 1 0 16500 0 1 15400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_525
timestamp 1675431769
transform 1 0 16500 0 1 16500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_526
timestamp 1675431769
transform 1 0 16500 0 1 17600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_527
timestamp 1675431769
transform 1 0 17050 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_528
timestamp 1675431769
transform 1 0 17050 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_529
timestamp 1675431769
transform 1 0 17050 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_530
timestamp 1675431769
transform 1 0 17050 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_531
timestamp 1675431769
transform 1 0 17050 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_532
timestamp 1675431769
transform 1 0 17050 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_533
timestamp 1675431769
transform 1 0 17050 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_534
timestamp 1675431769
transform 1 0 17050 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_535
timestamp 1675431769
transform 1 0 17050 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_536
timestamp 1675431769
transform 1 0 17050 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_537
timestamp 1675431769
transform 1 0 17050 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_538
timestamp 1675431769
transform 1 0 17050 0 1 12650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_539
timestamp 1675431769
transform 1 0 17050 0 1 13750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_540
timestamp 1675431769
transform 1 0 17050 0 1 14850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_541
timestamp 1675431769
transform 1 0 17050 0 1 15950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_542
timestamp 1675431769
transform 1 0 17050 0 1 17050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_543
timestamp 1675431769
transform 1 0 17050 0 1 18150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_544
timestamp 1675431769
transform 1 0 17600 0 1 0
box -113 -113 663 663
use nmos_source_in  nmos_source_in_545
timestamp 1675431769
transform 1 0 17600 0 1 1100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_546
timestamp 1675431769
transform 1 0 17600 0 1 2200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_547
timestamp 1675431769
transform 1 0 17600 0 1 3300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_548
timestamp 1675431769
transform 1 0 17600 0 1 4400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_549
timestamp 1675431769
transform 1 0 17600 0 1 5500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_550
timestamp 1675431769
transform 1 0 17600 0 1 6600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_551
timestamp 1675431769
transform 1 0 17600 0 1 7700
box -113 -113 663 663
use nmos_source_in  nmos_source_in_552
timestamp 1675431769
transform 1 0 17600 0 1 8800
box -113 -113 663 663
use nmos_source_in  nmos_source_in_553
timestamp 1675431769
transform 1 0 17600 0 1 9900
box -113 -113 663 663
use nmos_source_in  nmos_source_in_554
timestamp 1675431769
transform 1 0 17600 0 1 11000
box -113 -113 663 663
use nmos_source_in  nmos_source_in_555
timestamp 1675431769
transform 1 0 17600 0 1 12100
box -113 -113 663 663
use nmos_source_in  nmos_source_in_556
timestamp 1675431769
transform 1 0 17600 0 1 13200
box -113 -113 663 663
use nmos_source_in  nmos_source_in_557
timestamp 1675431769
transform 1 0 17600 0 1 14300
box -113 -113 663 663
use nmos_source_in  nmos_source_in_558
timestamp 1675431769
transform 1 0 17600 0 1 15400
box -113 -113 663 663
use nmos_source_in  nmos_source_in_559
timestamp 1675431769
transform 1 0 17600 0 1 16500
box -113 -113 663 663
use nmos_source_in  nmos_source_in_560
timestamp 1675431769
transform 1 0 17600 0 1 17600
box -113 -113 663 663
use nmos_source_in  nmos_source_in_561
timestamp 1675431769
transform 1 0 18150 0 1 550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_562
timestamp 1675431769
transform 1 0 18150 0 1 1650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_563
timestamp 1675431769
transform 1 0 18150 0 1 2750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_564
timestamp 1675431769
transform 1 0 18150 0 1 3850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_565
timestamp 1675431769
transform 1 0 18150 0 1 4950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_566
timestamp 1675431769
transform 1 0 18150 0 1 6050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_567
timestamp 1675431769
transform 1 0 18150 0 1 7150
box -113 -113 663 663
use nmos_source_in  nmos_source_in_568
timestamp 1675431769
transform 1 0 18150 0 1 8250
box -113 -113 663 663
use nmos_source_in  nmos_source_in_569
timestamp 1675431769
transform 1 0 18150 0 1 9350
box -113 -113 663 663
use nmos_source_in  nmos_source_in_570
timestamp 1675431769
transform 1 0 18150 0 1 10450
box -113 -113 663 663
use nmos_source_in  nmos_source_in_571
timestamp 1675431769
transform 1 0 18150 0 1 11550
box -113 -113 663 663
use nmos_source_in  nmos_source_in_572
timestamp 1675431769
transform 1 0 18150 0 1 12650
box -113 -113 663 663
use nmos_source_in  nmos_source_in_573
timestamp 1675431769
transform 1 0 18150 0 1 13750
box -113 -113 663 663
use nmos_source_in  nmos_source_in_574
timestamp 1675431769
transform 1 0 18150 0 1 14850
box -113 -113 663 663
use nmos_source_in  nmos_source_in_575
timestamp 1675431769
transform 1 0 18150 0 1 15950
box -113 -113 663 663
use nmos_source_in  nmos_source_in_576
timestamp 1675431769
transform 1 0 18150 0 1 17050
box -113 -113 663 663
use nmos_source_in  nmos_source_in_577
timestamp 1675431769
transform 1 0 18150 0 1 18150
box -113 -113 663 663
<< properties >>
string MASKHINTS_HVI -280 74800 0 75080 -280 -280 0 0 74800 -280 75080 0 74800 74800 75080 75080
string MASKHINTS_HVNTM -2014 -2214 -42 -2158 -2014 -2158 -1958 -242 75042 76758 77014 76814 76958 74842 77014 76758 -340 74860 -60 75140
<< end >>
