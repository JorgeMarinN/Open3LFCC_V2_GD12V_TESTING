magic
tech sky130A
timestamp 1698272741
<< mvnmos >>
rect 29 13 79 413
rect 108 13 158 413
rect 187 13 237 413
rect 266 13 316 413
rect 345 13 395 413
rect 424 13 474 413
rect 503 13 553 413
rect 582 13 632 413
rect 661 13 711 413
rect 740 13 790 413
rect 819 13 869 413
rect 898 13 948 413
rect 977 13 1027 413
rect 1056 13 1106 413
rect 1135 13 1185 413
rect 1214 13 1264 413
rect 1293 13 1343 413
rect 1372 13 1422 413
<< mvndiff >>
rect 0 407 29 413
rect 0 19 6 407
rect 23 19 29 407
rect 0 13 29 19
rect 79 407 108 413
rect 79 19 85 407
rect 102 19 108 407
rect 79 13 108 19
rect 158 407 187 413
rect 158 19 164 407
rect 181 19 187 407
rect 158 13 187 19
rect 237 407 266 413
rect 237 19 243 407
rect 260 19 266 407
rect 237 13 266 19
rect 316 407 345 413
rect 316 19 322 407
rect 339 19 345 407
rect 316 13 345 19
rect 395 407 424 413
rect 395 19 401 407
rect 418 19 424 407
rect 395 13 424 19
rect 474 407 503 413
rect 474 19 480 407
rect 497 19 503 407
rect 474 13 503 19
rect 553 407 582 413
rect 553 19 559 407
rect 576 19 582 407
rect 553 13 582 19
rect 632 407 661 413
rect 632 19 638 407
rect 655 19 661 407
rect 632 13 661 19
rect 711 407 740 413
rect 711 19 717 407
rect 734 19 740 407
rect 711 13 740 19
rect 790 407 819 413
rect 790 19 796 407
rect 813 19 819 407
rect 790 13 819 19
rect 869 407 898 413
rect 869 19 875 407
rect 892 19 898 407
rect 869 13 898 19
rect 948 407 977 413
rect 948 19 954 407
rect 971 19 977 407
rect 948 13 977 19
rect 1027 407 1056 413
rect 1027 19 1033 407
rect 1050 19 1056 407
rect 1027 13 1056 19
rect 1106 407 1135 413
rect 1106 19 1112 407
rect 1129 19 1135 407
rect 1106 13 1135 19
rect 1185 407 1214 413
rect 1185 19 1191 407
rect 1208 19 1214 407
rect 1185 13 1214 19
rect 1264 407 1293 413
rect 1264 19 1270 407
rect 1287 19 1293 407
rect 1264 13 1293 19
rect 1343 407 1372 413
rect 1343 19 1349 407
rect 1366 19 1372 407
rect 1343 13 1372 19
rect 1422 407 1451 413
rect 1422 19 1428 407
rect 1445 19 1451 407
rect 1422 13 1451 19
<< mvndiffc >>
rect 6 19 23 407
rect 85 19 102 407
rect 164 19 181 407
rect 243 19 260 407
rect 322 19 339 407
rect 401 19 418 407
rect 480 19 497 407
rect 559 19 576 407
rect 638 19 655 407
rect 717 19 734 407
rect 796 19 813 407
rect 875 19 892 407
rect 954 19 971 407
rect 1033 19 1050 407
rect 1112 19 1129 407
rect 1191 19 1208 407
rect 1270 19 1287 407
rect 1349 19 1366 407
rect 1428 19 1445 407
<< poly >>
rect 29 413 79 426
rect 108 413 158 426
rect 187 413 237 426
rect 266 413 316 426
rect 345 413 395 426
rect 424 413 474 426
rect 503 413 553 426
rect 582 413 632 426
rect 661 413 711 426
rect 740 413 790 426
rect 819 413 869 426
rect 898 413 948 426
rect 977 413 1027 426
rect 1056 413 1106 426
rect 1135 413 1185 426
rect 1214 413 1264 426
rect 1293 413 1343 426
rect 1372 413 1422 426
rect 29 0 79 13
rect 108 0 158 13
rect 187 0 237 13
rect 266 0 316 13
rect 345 0 395 13
rect 424 0 474 13
rect 503 0 553 13
rect 582 0 632 13
rect 661 0 711 13
rect 740 0 790 13
rect 819 0 869 13
rect 898 0 948 13
rect 977 0 1027 13
rect 1056 0 1106 13
rect 1135 0 1185 13
rect 1214 0 1264 13
rect 1293 0 1343 13
rect 1372 0 1422 13
<< locali >>
rect 6 407 23 415
rect 6 11 23 19
rect 85 407 102 415
rect 85 11 102 19
rect 164 407 181 415
rect 164 11 181 19
rect 243 407 260 415
rect 243 11 260 19
rect 322 407 339 415
rect 322 11 339 19
rect 401 407 418 415
rect 401 11 418 19
rect 480 407 497 415
rect 480 11 497 19
rect 559 407 576 415
rect 559 11 576 19
rect 638 407 655 415
rect 638 11 655 19
rect 717 407 734 415
rect 717 11 734 19
rect 796 407 813 415
rect 796 11 813 19
rect 875 407 892 415
rect 875 11 892 19
rect 954 407 971 415
rect 954 11 971 19
rect 1033 407 1050 415
rect 1033 11 1050 19
rect 1112 407 1129 415
rect 1112 11 1129 19
rect 1191 407 1208 415
rect 1191 11 1208 19
rect 1270 407 1287 415
rect 1270 11 1287 19
rect 1349 407 1366 415
rect 1349 11 1366 19
rect 1428 407 1445 415
rect 1428 11 1445 19
<< viali >>
rect 6 19 23 407
rect 85 19 102 407
rect 164 19 181 407
rect 243 19 260 407
rect 322 19 339 407
rect 401 19 418 407
rect 480 19 497 407
rect 559 19 576 407
rect 638 19 655 407
rect 717 19 734 407
rect 796 19 813 407
rect 875 19 892 407
rect 954 19 971 407
rect 1033 19 1050 407
rect 1112 19 1129 407
rect 1191 19 1208 407
rect 1270 19 1287 407
rect 1349 19 1366 407
rect 1428 19 1445 407
<< metal1 >>
rect 3 407 26 413
rect 3 19 6 407
rect 23 19 26 407
rect 3 13 26 19
rect 82 407 105 413
rect 82 19 85 407
rect 102 19 105 407
rect 82 13 105 19
rect 161 407 184 413
rect 161 19 164 407
rect 181 19 184 407
rect 161 13 184 19
rect 240 407 263 413
rect 240 19 243 407
rect 260 19 263 407
rect 240 13 263 19
rect 319 407 342 413
rect 319 19 322 407
rect 339 19 342 407
rect 319 13 342 19
rect 398 407 421 413
rect 398 19 401 407
rect 418 19 421 407
rect 398 13 421 19
rect 477 407 500 413
rect 477 19 480 407
rect 497 19 500 407
rect 477 13 500 19
rect 556 407 579 413
rect 556 19 559 407
rect 576 19 579 407
rect 556 13 579 19
rect 635 407 658 413
rect 635 19 638 407
rect 655 19 658 407
rect 635 13 658 19
rect 714 407 737 413
rect 714 19 717 407
rect 734 19 737 407
rect 714 13 737 19
rect 793 407 816 413
rect 793 19 796 407
rect 813 19 816 407
rect 793 13 816 19
rect 872 407 895 413
rect 872 19 875 407
rect 892 19 895 407
rect 872 13 895 19
rect 951 407 974 413
rect 951 19 954 407
rect 971 19 974 407
rect 951 13 974 19
rect 1030 407 1053 413
rect 1030 19 1033 407
rect 1050 19 1053 407
rect 1030 13 1053 19
rect 1109 407 1132 413
rect 1109 19 1112 407
rect 1129 19 1132 407
rect 1109 13 1132 19
rect 1188 407 1211 413
rect 1188 19 1191 407
rect 1208 19 1211 407
rect 1188 13 1211 19
rect 1267 407 1290 413
rect 1267 19 1270 407
rect 1287 19 1290 407
rect 1267 13 1290 19
rect 1346 407 1369 413
rect 1346 19 1349 407
rect 1366 19 1369 407
rect 1346 13 1369 19
rect 1425 407 1448 413
rect 1425 19 1428 407
rect 1445 19 1448 407
rect 1425 13 1448 19
<< end >>
