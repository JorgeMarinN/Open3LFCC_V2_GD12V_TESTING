magic
tech sky130A
magscale 1 2
timestamp 1700236551
<< checkpaint >>
rect -1037 1671 1512 2181
rect -1193 1557 1512 1671
rect -1193 -997 1546 1557
rect -1193 -1101 1361 -997
<< nwell >>
rect 0 309 5760 867
<< locali >>
rect 223 879 252 921
rect 5537 879 5846 921
rect 67 377 101 411
rect 5786 305 5846 879
rect 252 263 286 297
rect 5647 263 5846 305
rect 67 159 101 193
<< metal1 >>
rect -300 1088 38 1184
rect -300 96 -200 1088
rect -300 0 38 96
use sp_delay  sp_delay_0
timestamp 1700230441
transform 1 0 38 0 1 48
box -38 -48 5722 592
use sp_delay  sp_delay_1
timestamp 1700230441
transform -1 0 5722 0 -1 1136
box -38 -48 5722 592
<< labels >>
rlabel locali 67 377 101 411 5 VCC
port 1 s
rlabel locali 67 159 101 193 5 VSS
port 2 s
rlabel locali 252 263 286 297 5 VIN
port 3 s
rlabel locali 223 879 252 921 5 VOUT
port 4 s
<< end >>
