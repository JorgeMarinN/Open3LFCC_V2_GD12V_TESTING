magic
tech sky130A
timestamp 1698869965
<< mvnmos >>
rect -140 -129 160 371
rect 189 -129 489 371
<< mvndiff >>
rect -169 365 -140 371
rect -169 -123 -163 365
rect -146 -123 -140 365
rect -169 -129 -140 -123
rect 160 365 189 371
rect 160 -123 166 365
rect 183 -123 189 365
rect 160 -129 189 -123
rect 489 365 518 371
rect 489 -123 495 365
rect 512 -123 518 365
rect 489 -129 518 -123
<< mvndiffc >>
rect -163 -123 -146 365
rect 166 -123 183 365
rect 495 -123 512 365
<< poly >>
rect -140 371 160 384
rect 189 371 489 384
rect -140 -142 160 -129
rect 189 -142 489 -129
<< locali >>
rect -163 365 -146 373
rect -163 -131 -146 -123
rect 166 365 183 373
rect 166 -131 183 -123
rect 495 365 512 373
rect 495 -131 512 -123
<< viali >>
rect -163 -123 -146 365
rect 166 -123 183 365
rect 495 -123 512 365
<< metal1 >>
rect -166 365 -143 371
rect -166 -123 -163 365
rect -146 -123 -143 365
rect -166 -129 -143 -123
rect 163 365 186 371
rect 163 -123 166 365
rect 183 -123 186 365
rect 163 -129 186 -123
rect 492 365 515 371
rect 492 -123 495 365
rect 512 -123 515 365
rect 492 -129 515 -123
<< end >>
