magic
tech sky130A
timestamp 1698778120
<< mvnmos >>
rect 29 13 229 413
rect 258 13 458 413
rect 487 13 687 413
<< mvndiff >>
rect 0 407 29 413
rect 0 19 6 407
rect 23 19 29 407
rect 0 13 29 19
rect 229 407 258 413
rect 229 19 235 407
rect 252 19 258 407
rect 229 13 258 19
rect 458 407 487 413
rect 458 19 464 407
rect 481 19 487 407
rect 458 13 487 19
rect 687 407 716 413
rect 687 19 693 407
rect 710 19 716 407
rect 687 13 716 19
<< mvndiffc >>
rect 6 19 23 407
rect 235 19 252 407
rect 464 19 481 407
rect 693 19 710 407
<< poly >>
rect 29 413 229 426
rect 258 413 458 426
rect 487 413 687 426
rect 29 0 229 13
rect 258 0 458 13
rect 487 0 687 13
<< locali >>
rect 6 407 23 415
rect 6 11 23 19
rect 235 407 252 415
rect 235 11 252 19
rect 464 407 481 415
rect 464 11 481 19
rect 693 407 710 415
rect 693 11 710 19
<< viali >>
rect 6 19 23 407
rect 235 19 252 407
rect 464 19 481 407
rect 693 19 710 407
<< metal1 >>
rect 3 407 26 413
rect 3 19 6 407
rect 23 19 26 407
rect 3 13 26 19
rect 232 407 255 413
rect 232 19 235 407
rect 252 19 255 407
rect 232 13 255 19
rect 461 407 484 413
rect 461 19 464 407
rect 481 19 484 407
rect 461 13 484 19
rect 690 407 713 413
rect 690 19 693 407
rect 710 19 713 407
rect 690 13 713 19
<< end >>
