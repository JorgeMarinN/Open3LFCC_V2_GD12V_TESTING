magic
tech sky130A
magscale 1 2
timestamp 1700236959
<< checkpaint >>
rect -7032 4496 1732 8592
rect -7032 628 1832 4496
rect -6432 -3468 1832 628
<< dnwell >>
rect -187 -1532 7721 108
<< nwell >>
rect -267 -98 7801 2502
rect -267 -1326 19 -98
rect 7515 -1326 7801 -98
rect -267 -1612 7801 -1326
<< pwell >>
rect 19 -1326 7515 -98
<< mvnsubdiff >>
rect -187 -196 -107 -166
rect -187 -1296 -167 -196
rect -127 -1296 -107 -196
rect -187 -1326 -107 -1296
rect 7641 -196 7721 -166
rect 7641 -1296 7661 -196
rect 7701 -1296 7721 -196
rect 7641 -1326 7721 -1296
rect 19 -1472 7515 -1452
rect 19 -1512 49 -1472
rect 7485 -1512 7515 -1472
rect 19 -1532 7515 -1512
<< mvnsubdiffcont >>
rect -167 -1296 -127 -196
rect 7661 -1296 7701 -196
rect 49 -1512 7485 -1472
<< locali >>
rect -187 200 99 300
rect 7435 200 7721 300
rect -187 -196 -107 200
rect -187 -1296 -167 -196
rect -127 -1296 -107 -196
rect -187 -1326 -107 -1296
rect 7641 -196 7721 200
rect 7641 -1296 7661 -196
rect 7701 -1296 7721 -196
rect 7641 -1326 7721 -1296
rect 19 -1472 7515 -1452
rect 19 -1512 49 -1472
rect 7485 -1512 7515 -1472
rect 19 -1532 7515 -1512
<< viali >>
rect -167 -1296 -127 -196
rect 7661 -1296 7701 -196
rect 49 -1512 7485 -1472
<< metal1 >>
rect -3100 4640 -3000 4660
rect -3100 4580 -3080 4640
rect -3020 4580 -3000 4640
rect -3100 4560 -3000 4580
rect -2480 3460 -2380 3480
rect -2480 3400 -2460 3460
rect -2400 3400 -2380 3460
rect -2480 3380 -2380 3400
rect -3586 2400 7468 2600
rect -1200 2180 -800 2200
rect -1200 2020 -1180 2180
rect -820 2020 -800 2180
rect -1200 -89 -800 2020
rect 660 1460 1060 2400
rect 2500 1460 2900 2400
rect 66 1260 4340 1460
rect 1400 16 2200 116
rect 3200 96 3680 116
rect 3296 36 3680 96
rect 3200 16 3680 36
rect -1400 -1160 -800 -89
rect -634 -32 1140 -12
rect -634 -92 -614 -32
rect -554 -92 1140 -32
rect -634 -112 1140 -92
rect -207 -196 -107 -166
rect -207 -1296 -167 -196
rect -127 -1296 -107 -196
rect 1738 -1060 1838 16
rect 3580 -824 3680 16
rect 3580 -884 3600 -824
rect 3660 -884 3680 -824
rect 3580 -904 3680 -884
rect 7641 -196 7741 -166
rect 1738 -1120 1758 -1060
rect 1818 -1120 1838 -1060
rect 1738 -1140 1838 -1120
rect 3730 -1076 4320 -980
rect 3730 -1220 7488 -1076
rect -207 -1452 -107 -1296
rect 46 -1300 7488 -1220
rect 7641 -1296 7661 -196
rect 7701 -1296 7741 -196
rect 7641 -1452 7741 -1296
rect -207 -1472 7741 -1452
rect -207 -1512 49 -1472
rect 7485 -1512 7741 -1472
rect -207 -1552 7741 -1512
<< via1 >>
rect -3080 4580 -3020 4640
rect -2460 3400 -2400 3460
rect -1180 2820 -820 2876
rect -1180 2020 -820 2180
rect 280 36 796 96
rect 2780 36 3296 96
rect -614 -92 -554 -32
rect 2780 -92 3296 -32
rect 3600 -884 3660 -824
rect 1758 -1120 1818 -1060
<< metal2 >>
rect -3100 4640 -3000 4660
rect -3100 4580 -3080 4640
rect -3020 4580 -3000 4640
rect -3100 4560 -3000 4580
rect -2480 3460 -2380 3480
rect -2480 3400 -2460 3460
rect -2400 3400 -2380 3460
rect -2480 3380 -2380 3400
rect -1200 2876 -800 2896
rect -1200 2820 -1180 2876
rect -820 2820 -800 2876
rect -1200 2180 -800 2820
rect -1200 2020 -1180 2180
rect -820 2020 -800 2180
rect -1200 2000 -800 2020
rect -1734 1118 -394 1218
rect -1734 990 -534 1090
rect -634 -32 -534 990
rect -634 -92 -614 -32
rect -554 -92 -534 -32
rect -634 -112 -534 -92
rect -494 -12 -394 1118
rect 260 96 3316 116
rect 260 36 280 96
rect 796 36 2780 96
rect 3296 36 3316 96
rect 260 16 3316 36
rect -494 -32 3316 -12
rect -494 -92 2780 -32
rect 3296 -92 3316 -32
rect -494 -112 3316 -92
rect 3580 -824 4000 -804
rect 3580 -884 3600 -824
rect 3660 -884 4000 -824
rect 3580 -904 4000 -884
rect 1738 -1060 1838 -1040
rect 1738 -1120 1758 -1060
rect 1818 -1120 1838 -1060
rect 1738 -1300 1838 -1120
rect 4102 -1300 4202 -804
rect 1738 -1400 4202 -1300
<< via2 >>
rect -3080 4580 -3020 4640
rect -2460 3400 -2400 3460
rect -3280 484 -2920 544
rect -2480 484 -2120 544
<< metal3 >>
rect -3100 4640 -2200 4660
rect -3100 4580 -3080 4640
rect -3020 4580 -2200 4640
rect -3100 4560 -2200 4580
rect -3000 3460 -2380 3480
rect -3000 3400 -2460 3460
rect -2400 3400 -2380 3460
rect -3000 3380 -2380 3400
rect -3000 564 -2900 3380
rect -2300 564 -2200 4560
rect -3300 544 -2900 564
rect -3300 484 -3280 544
rect -2920 484 -2900 544
rect -3300 464 -2900 484
rect -2500 544 -2100 564
rect -2500 484 -2480 544
rect -2120 484 -2100 544
rect -2500 464 -2100 484
use boot_ls_stage  boot_ls_stage_0
timestamp 1699931927
transform 1 0 -2811 0 1 1104
box -1778 -2264 1444 1422
use buffer  buffer_0
timestamp 1699046184
transform 1 0 4051 0 1 -12
box -395 -1088 3503 2502
use nand_5v  nand_5v_0
timestamp 1699971027
transform 1 0 867 0 1 2
box -867 -1302 867 1348
use nand_5v  nand_5v_1
timestamp 1699971027
transform 1 0 2709 0 1 2
box -867 -1302 867 1348
use short_pulse_generator  short_pulse_generator_0
timestamp 1700236738
transform 0 -1 -2200 -1 0 6160
box -38 -6380 3360 1140
<< labels >>
rlabel metal1 7200 -1300 7400 -1100 5 VSource
rlabel metal1 -3586 2400 -3386 2600 1 VBOOT
<< end >>
