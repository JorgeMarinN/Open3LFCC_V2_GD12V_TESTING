magic
tech sky130A
magscale 1 2
timestamp 1699928925
<< xpolycontact >>
rect -60 1040 10 1472
rect -60 86 10 518
rect 106 1040 176 1472
rect 106 86 176 518
rect 272 1040 342 1472
rect 272 86 342 518
rect 438 1040 508 1472
rect 438 86 508 518
rect 604 1040 674 1472
rect 604 86 674 518
<< xpolyres >>
rect -60 518 10 1040
rect 106 518 176 1040
rect 272 518 342 1040
rect 438 518 508 1040
rect 604 518 674 1040
<< viali >>
rect -44 1057 -6 1454
rect 122 1057 160 1454
rect 288 1057 326 1454
rect 454 1057 492 1454
rect 620 1057 658 1454
rect -44 104 -6 501
rect 122 104 160 501
rect 288 104 326 501
rect 454 104 492 501
rect 620 104 658 501
<< metal1 >>
rect -50 1454 0 1466
rect -50 1057 -44 1454
rect -6 1057 0 1454
rect -50 1045 0 1057
rect 116 1454 166 1466
rect 116 1057 122 1454
rect 160 1057 166 1454
rect 116 1045 166 1057
rect 282 1454 332 1466
rect 282 1057 288 1454
rect 326 1057 332 1454
rect 282 1045 332 1057
rect 448 1454 498 1466
rect 448 1057 454 1454
rect 492 1057 498 1454
rect 448 1045 498 1057
rect 614 1454 664 1466
rect 614 1057 620 1454
rect 658 1057 664 1454
rect 614 1045 664 1057
rect -50 501 0 513
rect -50 104 -44 501
rect -6 104 0 501
rect -50 92 0 104
rect 116 501 166 513
rect 116 104 122 501
rect 160 104 166 501
rect 116 92 166 104
rect 282 501 332 513
rect 282 104 288 501
rect 326 104 332 501
rect 282 92 332 104
rect 448 501 498 513
rect 448 104 454 501
rect 492 104 498 501
rect 448 92 498 104
rect 614 501 664 513
rect 614 104 620 501
rect 658 104 664 501
rect 614 92 664 104
<< res0p35 >>
rect -62 516 12 1042
rect 104 516 178 1042
rect 270 516 344 1042
rect 436 516 510 1042
rect 602 516 676 1042
<< end >>
