magic
tech sky130A
timestamp 1698625803
<< nwell >>
rect -117 -61 1268 105
<< mvpmos >>
rect -55 -28 45 72
rect 74 -28 174 72
rect 203 -28 303 72
rect 332 -28 432 72
rect 461 -28 561 72
rect 590 -28 690 72
rect 719 -28 819 72
rect 848 -28 948 72
rect 977 -28 1077 72
rect 1106 -28 1206 72
<< mvpdiff >>
rect -84 66 -55 72
rect -84 -22 -78 66
rect -61 -22 -55 66
rect -84 -28 -55 -22
rect 45 66 74 72
rect 45 -22 51 66
rect 68 -22 74 66
rect 45 -28 74 -22
rect 174 66 203 72
rect 174 -22 180 66
rect 197 -22 203 66
rect 174 -28 203 -22
rect 303 66 332 72
rect 303 -22 309 66
rect 326 -22 332 66
rect 303 -28 332 -22
rect 432 66 461 72
rect 432 -22 438 66
rect 455 -22 461 66
rect 432 -28 461 -22
rect 561 66 590 72
rect 561 -22 567 66
rect 584 -22 590 66
rect 561 -28 590 -22
rect 690 66 719 72
rect 690 -22 696 66
rect 713 -22 719 66
rect 690 -28 719 -22
rect 819 66 848 72
rect 819 -22 825 66
rect 842 -22 848 66
rect 819 -28 848 -22
rect 948 66 977 72
rect 948 -22 954 66
rect 971 -22 977 66
rect 948 -28 977 -22
rect 1077 66 1106 72
rect 1077 -22 1083 66
rect 1100 -22 1106 66
rect 1077 -28 1106 -22
rect 1206 66 1235 72
rect 1206 -22 1212 66
rect 1229 -22 1235 66
rect 1206 -28 1235 -22
<< mvpdiffc >>
rect -78 -22 -61 66
rect 51 -22 68 66
rect 180 -22 197 66
rect 309 -22 326 66
rect 438 -22 455 66
rect 567 -22 584 66
rect 696 -22 713 66
rect 825 -22 842 66
rect 954 -22 971 66
rect 1083 -22 1100 66
rect 1212 -22 1229 66
<< poly >>
rect -55 72 45 85
rect 74 72 174 85
rect 203 72 303 85
rect 332 72 432 85
rect 461 72 561 85
rect 590 72 690 85
rect 719 72 819 85
rect 848 72 948 85
rect 977 72 1077 85
rect 1106 72 1206 85
rect -55 -41 45 -28
rect 74 -41 174 -28
rect 203 -41 303 -28
rect 332 -41 432 -28
rect 461 -41 561 -28
rect 590 -41 690 -28
rect 719 -41 819 -28
rect 848 -41 948 -28
rect 977 -41 1077 -28
rect 1106 -41 1206 -28
<< locali >>
rect -78 66 -61 74
rect -78 -30 -61 -22
rect 51 66 68 74
rect 51 -30 68 -22
rect 180 66 197 74
rect 180 -30 197 -22
rect 309 66 326 74
rect 309 -30 326 -22
rect 438 66 455 74
rect 438 -30 455 -22
rect 567 66 584 74
rect 567 -30 584 -22
rect 696 66 713 74
rect 696 -30 713 -22
rect 825 66 842 74
rect 825 -30 842 -22
rect 954 66 971 74
rect 954 -30 971 -22
rect 1083 66 1100 74
rect 1083 -30 1100 -22
rect 1212 66 1229 74
rect 1212 -30 1229 -22
<< viali >>
rect -78 -22 -61 66
rect 51 -22 68 66
rect 180 -22 197 66
rect 309 -22 326 66
rect 438 -22 455 66
rect 567 -22 584 66
rect 696 -22 713 66
rect 825 -22 842 66
rect 954 -22 971 66
rect 1083 -22 1100 66
rect 1212 -22 1229 66
<< metal1 >>
rect -81 66 -58 72
rect -81 -22 -78 66
rect -61 -22 -58 66
rect -81 -28 -58 -22
rect 48 66 71 72
rect 48 -22 51 66
rect 68 -22 71 66
rect 48 -28 71 -22
rect 177 66 200 72
rect 177 -22 180 66
rect 197 -22 200 66
rect 177 -28 200 -22
rect 306 66 329 72
rect 306 -22 309 66
rect 326 -22 329 66
rect 306 -28 329 -22
rect 435 66 458 72
rect 435 -22 438 66
rect 455 -22 458 66
rect 435 -28 458 -22
rect 564 66 587 72
rect 564 -22 567 66
rect 584 -22 587 66
rect 564 -28 587 -22
rect 693 66 716 72
rect 693 -22 696 66
rect 713 -22 716 66
rect 693 -28 716 -22
rect 822 66 845 72
rect 822 -22 825 66
rect 842 -22 845 66
rect 822 -28 845 -22
rect 951 66 974 72
rect 951 -22 954 66
rect 971 -22 974 66
rect 951 -28 974 -22
rect 1080 66 1103 72
rect 1080 -22 1083 66
rect 1100 -22 1103 66
rect 1080 -28 1103 -22
rect 1209 66 1232 72
rect 1209 -22 1212 66
rect 1229 -22 1232 66
rect 1209 -28 1232 -22
<< end >>
