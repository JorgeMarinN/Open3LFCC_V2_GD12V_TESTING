magic
tech sky130A
timestamp 1698627441
<< nwell >>
rect -30 -4 581 312
<< mvpmos >>
rect 32 29 132 279
rect 161 29 261 279
rect 290 29 390 279
rect 419 29 519 279
<< mvpdiff >>
rect 3 273 32 279
rect 3 35 9 273
rect 26 35 32 273
rect 3 29 32 35
rect 132 273 161 279
rect 132 35 138 273
rect 155 35 161 273
rect 132 29 161 35
rect 261 273 290 279
rect 261 35 267 273
rect 284 35 290 273
rect 261 29 290 35
rect 390 273 419 279
rect 390 35 396 273
rect 413 35 419 273
rect 390 29 419 35
rect 519 273 548 279
rect 519 35 525 273
rect 542 35 548 273
rect 519 29 548 35
<< mvpdiffc >>
rect 9 35 26 273
rect 138 35 155 273
rect 267 35 284 273
rect 396 35 413 273
rect 525 35 542 273
<< poly >>
rect 32 279 132 292
rect 161 279 261 292
rect 290 279 390 292
rect 419 279 519 292
rect 32 16 132 29
rect 161 16 261 29
rect 290 16 390 29
rect 419 16 519 29
<< locali >>
rect 9 273 26 281
rect 9 27 26 35
rect 138 273 155 281
rect 138 27 155 35
rect 267 273 284 281
rect 267 27 284 35
rect 396 273 413 281
rect 396 27 413 35
rect 525 273 542 281
rect 525 27 542 35
<< viali >>
rect 9 35 26 273
rect 138 35 155 273
rect 267 35 284 273
rect 396 35 413 273
rect 525 35 542 273
<< metal1 >>
rect 6 273 29 279
rect 6 35 9 273
rect 26 35 29 273
rect 6 29 29 35
rect 135 273 158 279
rect 135 35 138 273
rect 155 35 158 273
rect 135 29 158 35
rect 264 273 287 279
rect 264 35 267 273
rect 284 35 287 273
rect 264 29 287 35
rect 393 273 416 279
rect 393 35 396 273
rect 413 35 416 273
rect 393 29 416 35
rect 522 273 545 279
rect 522 35 525 273
rect 542 35 545 273
rect 522 29 545 35
<< end >>
