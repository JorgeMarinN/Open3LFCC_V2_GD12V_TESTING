magic
tech sky130A
magscale 1 2
timestamp 1700237874
<< obsactive >>
rect -18000 61200 141200 79200
rect -18000 -18000 0 61200
rect 123200 -18000 141200 61200
<< metal1 >>
rect 6000 -620 6320 -600
rect 6000 -4080 6020 -620
rect 6000 -4200 6320 -4080
rect 15008 -620 15400 -600
rect 15008 -6420 15020 -620
rect 15380 -6420 15400 -620
rect 111200 -4620 111500 -4600
rect 111200 -4780 111220 -4620
rect 111480 -4780 111500 -4620
rect 111200 -4800 111500 -4780
rect 15008 -6600 15400 -6420
rect 4000 -6820 9600 -6800
rect 4000 -7180 9220 -6820
rect 9580 -7180 9600 -6820
rect 4000 -7200 9600 -7180
rect 111600 -10020 112000 -10000
rect 111600 -12800 111620 -10020
rect 111980 -12800 112000 -10020
rect 111600 -12824 112000 -12800
rect 112220 -12800 112320 -12780
rect 112220 -13200 112240 -12800
rect 112300 -13200 112320 -12800
rect 112220 -13220 112320 -13200
rect 9200 -44820 117000 -44800
rect 9200 -45180 9220 -44820
rect 9580 -45180 116620 -44820
rect 116980 -45180 117000 -44820
rect 9200 -45200 117000 -45180
rect 5800 -45420 112000 -45400
rect 5800 -45980 5820 -45420
rect 6380 -45980 111620 -45420
rect 111980 -45980 112000 -45420
rect 5800 -46000 112000 -45980
rect 15000 -46220 116000 -46200
rect 15000 -47180 15020 -46220
rect 15380 -47180 112220 -46220
rect 112380 -47180 116000 -46220
rect 15000 -47200 116000 -47180
<< via1 >>
rect 6020 -4080 6320 -620
rect 9400 -6000 9454 -5500
rect 15020 -6420 15380 -620
rect 111740 -4180 111980 -1160
rect 111220 -4780 111480 -4620
rect 9220 -7180 9580 -6820
rect 115432 -9280 115592 -8920
rect 111620 -12800 111980 -10020
rect 116620 -11403 116980 -11347
rect 112240 -13200 112300 -12800
rect 112220 -17200 112374 -14220
rect 112640 -16760 114760 -14640
rect 9220 -45180 9580 -44820
rect 116620 -45180 116980 -44820
rect 5820 -45980 6380 -45420
rect 111620 -45980 111980 -45420
rect 15020 -47180 15380 -46220
rect 112220 -47180 112380 -46220
<< metal2 >>
rect 58000 56000 66000 60000
rect 113000 6560 113200 6600
rect 10434 6360 10754 6400
rect 10434 5440 10474 6360
rect 10714 5440 10754 6360
rect 113000 6040 113040 6560
rect 113160 6040 113200 6560
rect 5800 580 6400 600
rect 5800 20 5820 580
rect 6380 20 6400 580
rect 5800 -620 6400 20
rect 5800 -4080 6020 -620
rect 6320 -4080 6400 -620
rect 10434 -800 10754 5440
rect 58000 2000 66000 6000
rect 111600 580 112000 600
rect 111600 40 111640 580
rect 111960 40 112000 580
rect 15000 -620 15400 -600
rect 5800 -45420 6400 -4080
rect 9384 -6000 9400 -5500
rect 9454 -6000 9470 -5500
rect 9384 -6800 9470 -6000
rect 15000 -6420 15020 -620
rect 15380 -6420 15400 -620
rect 111600 -1160 112000 40
rect 111600 -4180 111740 -1160
rect 111980 -4180 112000 -1160
rect 113000 -1200 113200 6040
rect 111600 -4200 112000 -4180
rect 111200 -4620 111500 -4600
rect 111200 -4780 111220 -4620
rect 111480 -4780 111500 -4620
rect 111200 -4800 111500 -4780
rect 9200 -6820 9600 -6800
rect 9200 -7180 9220 -6820
rect 9580 -7180 9600 -6820
rect 9200 -44820 9600 -7180
rect 9200 -45180 9220 -44820
rect 9580 -45180 9600 -44820
rect 9200 -45200 9600 -45180
rect 5800 -45980 5820 -45420
rect 6380 -45980 6400 -45420
rect 5800 -46000 6400 -45980
rect 15000 -46220 15400 -6420
rect 115412 -8920 115612 -8900
rect 115412 -9280 115432 -8920
rect 115592 -9280 115612 -8920
rect 115412 -9300 115612 -9280
rect 111600 -10020 112000 -10000
rect 111600 -12800 111620 -10020
rect 111980 -12800 112000 -10020
rect 116600 -11347 117000 -11327
rect 116600 -11403 116620 -11347
rect 116980 -11403 117000 -11347
rect 111600 -45420 112000 -12800
rect 112220 -12800 112320 -12780
rect 112220 -13200 112240 -12800
rect 112300 -13200 112320 -12800
rect 112220 -14200 112320 -13200
rect 111600 -45980 111620 -45420
rect 111980 -45980 112000 -45420
rect 111600 -46000 112000 -45980
rect 112200 -14220 112400 -14200
rect 112200 -17200 112220 -14220
rect 112374 -17200 112400 -14220
rect 112600 -14640 114800 -14600
rect 112600 -16760 112640 -14640
rect 114760 -16760 114800 -14640
rect 112600 -16800 114800 -16760
rect 15000 -47180 15020 -46220
rect 15380 -47180 15400 -46220
rect 15000 -47200 15400 -47180
rect 112200 -46220 112400 -17200
rect 116600 -44820 117000 -11403
rect 116600 -45180 116620 -44820
rect 116980 -45180 117000 -44820
rect 116600 -45200 117000 -45180
rect 112200 -47180 112220 -46220
rect 112380 -47180 112400 -46220
rect 112200 -47200 112400 -47180
<< via2 >>
rect 116000 54000 120000 58000
rect 10474 5440 10714 6360
rect 113040 6040 113160 6560
rect 5820 20 6380 580
rect 111640 40 111960 580
rect 113034 -3994 113094 -1462
rect 111220 -4780 111480 -4620
rect 115432 -9280 115592 -8920
rect 112640 -16760 114760 -14640
<< metal3 >>
rect 5800 580 6400 12000
rect 5800 20 5820 580
rect 6380 20 6400 580
rect 5800 0 6400 20
rect 10434 6360 10754 6400
rect 10434 5440 10474 6360
rect 10714 5440 10754 6360
rect 10434 -800 10754 5440
rect 22000 1560 108000 1600
rect 22000 440 22040 1560
rect 107960 440 108000 1560
rect 22000 0 108000 440
rect 111600 580 112000 6800
rect 111600 40 111640 580
rect 111960 40 112000 580
rect 111600 0 112000 40
rect 113000 6560 113200 6600
rect 113000 6040 113040 6560
rect 113160 6040 113200 6560
rect 113000 -1200 113200 6040
rect 113014 -1462 113114 -1200
rect 110000 -2040 111400 -2000
rect 110000 -43960 110040 -2040
rect 111360 -4600 111400 -2040
rect 113014 -3994 113034 -1462
rect 113094 -3994 113114 -1462
rect 113014 -4016 113114 -3994
rect 111360 -4620 111500 -4600
rect 111480 -4780 111500 -4620
rect 111360 -4800 111500 -4780
rect 111360 -8900 111400 -4800
rect 111360 -8920 115612 -8900
rect 111360 -9280 115432 -8920
rect 115592 -9280 115612 -8920
rect 111360 -9300 115612 -9280
rect 111360 -14600 111400 -9300
rect 111360 -14640 114800 -14600
rect 111360 -16760 112640 -14640
rect 114760 -16760 114800 -14640
rect 111360 -16800 114800 -16760
rect 111360 -43960 111400 -16800
rect 110000 -44000 111400 -43960
<< via3 >>
rect 116000 54000 120000 58000
rect 10474 5440 10714 6360
rect 22040 440 107960 1560
rect 110040 -4620 111360 -2040
rect 110040 -4780 111220 -4620
rect 111220 -4780 111360 -4620
rect 110040 -43960 111360 -4780
<< metal4 >>
rect 10434 6360 10754 6400
rect 10434 5440 10474 6360
rect 10714 5440 10754 6360
rect 10434 -800 10754 5440
rect 22000 1560 108000 2000
rect 22000 440 22040 1560
rect 107960 440 108000 1560
rect 22000 400 108000 440
rect 109320 -2040 111400 -2000
rect 109320 -43960 110040 -2040
rect 111360 -43960 111400 -2040
rect 109320 -44000 111400 -43960
<< via4 >>
rect 116000 54000 120000 58000
rect 10474 5440 10714 6360
rect 22040 440 107960 1560
<< metal5 >>
rect 2000 56000 6000 60000
rect 60000 46000 64000 50000
rect 10434 6360 10754 6400
rect 10434 5440 10474 6360
rect 10714 5440 10754 6360
rect 10434 -800 10754 5440
rect 22000 1560 108000 1600
rect 22000 440 22040 1560
rect 107960 440 108000 1560
rect 22000 0 108000 440
use bootstrap_diode  bootstrap_diode_0
timestamp 1700061388
transform -1 0 115130 0 1 -17114
box -286 -286 3102 3102
use driver_bootstrap  driver_bootstrap_0
timestamp 1700237389
transform 0 1 113012 1 0 -8631
box -4589 -1612 7801 6198
use level_shifter  level_shifter_0
timestamp 1666543010
transform 0 1 6200 1 0 -6600
box 0 0 6050 8936
use mimcap_210x420  mimcap_210x420_0
timestamp 1698868607
transform 1 0 20000 0 1 -44660
box 0 0 89320 44660
use power_stage_3  power_stage_3_0
timestamp 1699898483
transform 0 1 0 1 0 0
box 0 0 61200 123200
<< labels >>
rlabel metal5 2000 56000 6000 60000 1 VSS
rlabel metal5 116000 54000 120000 58000 1 VDD
rlabel metal5 60000 46000 64000 50000 1 Vout
rlabel metal1 4000 -7200 4400 -6800 7 V1v8
rlabel metal3 110000 -3400 111400 -2000 1 Vboot
rlabel metal1 115000 -47200 116000 -46200 3 V5v0LS
<< end >>
