magic
tech sky130A
timestamp 1700061388
<< dnwell >>
rect -103 -103 1511 1511
<< nwell >>
rect -143 1408 1551 1551
rect -143 0 0 1408
rect 1408 0 1551 1408
rect -143 -143 1551 0
<< pwell >>
rect 0 0 1408 1408
<< psubdiff >>
rect 18 1373 66 1390
rect 1342 1373 1390 1390
rect 18 35 35 1373
rect 1373 1342 1390 1373
rect 1373 35 1390 66
rect 18 18 66 35
rect 1342 18 1390 35
<< nsubdiff >>
rect 0 1435 15 1455
rect 1393 1435 1408 1455
rect 1435 1393 1455 1408
rect 1435 0 1455 15
rect 0 -47 15 -27
rect 1393 -47 1408 -27
<< psubdiffcont >>
rect 66 1373 1342 1390
rect 1373 66 1390 1342
rect 66 18 1342 35
<< nsubdiffcont >>
rect 15 1435 1393 1455
rect 1435 15 1455 1393
rect 15 -47 1393 -27
<< ndiode >>
rect 69 1333 1339 1339
rect 69 75 75 1333
rect 1333 75 1339 1333
rect 69 69 1339 75
<< ndiodec >>
rect 75 75 1333 1333
<< locali >>
rect 0 1435 15 1455
rect 1393 1435 1408 1455
rect 1435 1393 1455 1408
rect 18 1373 66 1390
rect 1342 1373 1390 1390
rect 18 35 35 1373
rect 1373 1342 1390 1373
rect 67 75 75 1333
rect 1333 75 1341 1333
rect 1373 35 1390 66
rect 18 18 66 35
rect 1342 18 1390 35
rect 1435 0 1455 15
rect 0 -47 15 -27
rect 1393 -47 1408 -27
<< viali >>
rect 15 1435 1393 1455
rect 66 1390 1342 1391
rect 66 1373 1342 1390
rect 75 75 1333 1333
rect 1373 66 1390 1342
rect 1390 66 1391 1342
rect 66 18 1342 35
rect 66 17 1342 18
rect 1435 15 1455 1393
rect 15 -47 1393 -27
<< metal1 >>
rect 0 1455 1465 1465
rect 0 1435 15 1455
rect 1393 1435 1465 1455
rect 0 1393 1465 1435
rect 0 1391 1435 1393
rect 0 1373 66 1391
rect 1342 1373 1435 1391
rect 0 1368 1435 1373
rect 1368 1342 1435 1368
rect 69 1333 1339 1336
rect 69 75 75 1333
rect 1333 75 1339 1333
rect 69 72 1339 75
rect 1368 66 1373 1342
rect 1391 66 1435 1342
rect 1368 40 1435 66
rect 0 35 1435 40
rect 0 17 66 35
rect 1342 17 1435 35
rect 0 15 1435 17
rect 1455 15 1465 1393
rect 0 -27 1465 15
rect 0 -47 15 -27
rect 1393 -47 1465 -27
rect 0 -57 1465 -47
<< end >>
