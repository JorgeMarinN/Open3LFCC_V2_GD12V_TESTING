magic
tech sky130A
timestamp 1699931197
<< viali >>
rect 474 463 491 481
rect 311 421 341 443
rect 428 426 446 443
rect 474 426 491 444
rect 903 429 921 447
rect 945 429 963 447
rect 996 429 1013 446
rect 94 63 113 137
rect 282 124 299 142
rect 1348 127 1365 145
rect 233 92 250 109
rect 281 81 298 99
rect 386 92 403 110
rect 477 92 495 109
rect 524 92 542 109
rect 569 92 587 109
rect 615 92 633 109
rect 661 93 679 110
rect 706 93 724 110
rect 754 92 771 110
rect 830 90 850 110
rect 923 92 942 109
rect 969 92 988 109
rect 1014 92 1033 109
rect 1060 92 1079 109
rect 1105 92 1124 109
rect 1148 92 1167 109
rect 1198 90 1217 110
rect 1301 90 1318 108
rect 1349 90 1366 108
rect 1448 90 1465 107
rect 1491 89 1508 106
rect 1538 88 1562 108
<< metal1 >>
rect 468 481 496 488
rect 468 463 474 481
rect 491 463 496 481
rect 468 454 496 463
rect 302 443 454 449
rect 302 421 311 443
rect 341 426 428 443
rect 446 426 454 443
rect 341 421 454 426
rect 302 414 454 421
rect 468 447 969 454
rect 468 444 903 447
rect 468 426 474 444
rect 491 429 903 444
rect 921 429 945 447
rect 963 429 969 447
rect 491 426 969 429
rect 468 424 969 426
rect 987 452 1024 454
rect 987 426 990 452
rect 1018 426 1024 452
rect 468 419 496 424
rect 987 420 1024 426
rect 1191 191 1231 192
rect 821 186 1231 191
rect 821 160 938 186
rect 966 160 989 186
rect 1017 160 1042 186
rect 1070 160 1231 186
rect 821 155 1231 160
rect 82 137 124 146
rect 82 63 94 137
rect 113 119 124 137
rect 276 142 349 148
rect 276 124 282 142
rect 299 135 349 142
rect 299 124 310 135
rect 113 109 258 119
rect 113 92 233 109
rect 250 92 258 109
rect 113 80 258 92
rect 276 99 310 124
rect 276 81 281 99
rect 298 92 310 99
rect 340 92 349 135
rect 298 81 349 92
rect 113 63 124 80
rect 276 76 349 81
rect 379 110 412 122
rect 379 92 386 110
rect 403 92 412 110
rect 276 75 304 76
rect 82 52 124 63
rect 379 56 412 92
rect 463 110 730 120
rect 463 109 661 110
rect 463 92 477 109
rect 495 92 524 109
rect 542 92 569 109
rect 587 92 615 109
rect 633 93 661 109
rect 679 93 706 110
rect 724 93 730 110
rect 633 92 730 93
rect 463 80 730 92
rect 744 110 777 125
rect 744 92 754 110
rect 771 92 777 110
rect 744 58 777 92
rect 821 110 861 155
rect 821 90 830 110
rect 850 90 861 110
rect 821 81 861 90
rect 912 114 1171 116
rect 912 109 1172 114
rect 912 92 923 109
rect 942 92 969 109
rect 988 92 1014 109
rect 1033 92 1060 109
rect 1079 92 1105 109
rect 1124 92 1148 109
rect 1167 92 1172 109
rect 912 85 1172 92
rect 1191 110 1231 155
rect 1191 90 1198 110
rect 1217 90 1231 110
rect 964 58 1087 85
rect 1191 82 1231 90
rect 1289 188 1327 192
rect 1289 161 1295 188
rect 1322 161 1327 188
rect 1289 108 1327 161
rect 1289 90 1301 108
rect 1318 90 1327 108
rect 1289 80 1327 90
rect 1342 145 1371 150
rect 1342 127 1348 145
rect 1365 129 1371 145
rect 1365 127 1514 129
rect 1342 108 1514 127
rect 1342 90 1349 108
rect 1366 107 1514 108
rect 1366 103 1448 107
rect 1366 90 1371 103
rect 1342 82 1371 90
rect 1437 90 1448 103
rect 1465 106 1514 107
rect 1465 90 1491 106
rect 1437 89 1491 90
rect 1508 89 1514 106
rect 1437 85 1514 89
rect 1530 108 1568 115
rect 1530 88 1538 108
rect 1562 88 1568 108
rect 1530 79 1568 88
rect 744 56 1179 58
rect 379 34 1179 56
rect 410 33 1179 34
rect 775 32 1179 33
<< rmetal1 >>
rect 1534 78 1568 79
<< via1 >>
rect 990 446 1018 452
rect 990 429 996 446
rect 996 429 1013 446
rect 1013 429 1018 446
rect 990 426 1018 429
rect 938 160 966 186
rect 989 160 1017 186
rect 1042 160 1070 186
rect 310 92 340 135
rect 1295 161 1322 188
<< metal2 >>
rect 982 452 1027 463
rect 303 135 349 449
rect 982 426 990 452
rect 1018 426 1027 452
rect 982 191 1027 426
rect 1090 191 1333 192
rect 926 188 1333 191
rect 926 186 1295 188
rect 926 160 938 186
rect 966 160 989 186
rect 1017 160 1042 186
rect 1070 161 1295 186
rect 1322 161 1333 188
rect 1070 160 1333 161
rect 926 157 1333 160
rect 926 156 1093 157
rect 303 92 310 135
rect 340 122 349 135
rect 340 120 738 122
rect 340 92 1574 120
rect 303 77 1574 92
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 889 0 1 319
box -19 -24 295 296
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_1
timestamp 1693170804
transform 1 0 1434 0 1 -21
box -19 -24 295 296
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 197 0 1 -19
box -19 -24 157 296
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1693170804
transform 1 0 389 0 1 316
box -19 -24 157 296
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1693170804
transform 1 0 1265 0 1 -20
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 29 0 1 -19
box -19 -24 157 296
use sky130_fd_sc_hd__inv_8  sky130_fd_sc_hd__inv_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 371 0 1 -18
box -19 -24 433 296
use sky130_fd_sc_hd__inv_8  sky130_fd_sc_hd__inv_8_1
timestamp 1693170804
transform 1 0 817 0 1 -19
box -19 -24 433 296
<< labels >>
rlabel space 1084 351 1110 553 1 VFE
rlabel space 1629 16 1655 218 1 VRE
rlabel space 38 87 69 114 1 VIN
<< end >>
