magic
tech sky130A
magscale 1 2
timestamp 1699971027
<< nwell >>
rect -867 102 867 1348
<< mvnmos >>
rect -629 -1168 -29 -168
rect 29 -1168 629 -168
<< mvpmos >>
rect -629 168 -29 1168
rect 29 168 629 1168
<< mvndiff >>
rect -687 -180 -629 -168
rect -687 -1156 -675 -180
rect -641 -1156 -629 -180
rect -687 -1168 -629 -1156
rect -29 -180 29 -168
rect -29 -1156 -17 -180
rect 17 -1156 29 -180
rect -29 -1168 29 -1156
rect 629 -180 687 -168
rect 629 -1156 641 -180
rect 675 -1156 687 -180
rect 629 -1168 687 -1156
<< mvpdiff >>
rect -687 1156 -629 1168
rect -687 180 -675 1156
rect -641 180 -629 1156
rect -687 168 -629 180
rect -29 1156 29 1168
rect -29 180 -17 1156
rect 17 180 29 1156
rect -29 168 29 180
rect 629 1156 687 1168
rect 629 180 641 1156
rect 675 180 687 1156
rect 629 168 687 180
<< mvndiffc >>
rect -675 -1156 -641 -180
rect -17 -1156 17 -180
rect 641 -1156 675 -180
<< mvpdiffc >>
rect -675 180 -641 1156
rect -17 180 17 1156
rect 641 180 675 1156
<< mvpsubdiff >>
rect -801 -198 -761 -168
rect -801 -1168 -761 -1138
rect 761 -198 801 -168
rect 761 -1168 801 -1138
rect -687 -1282 -657 -1242
rect 657 -1282 687 -1242
<< mvnsubdiff >>
rect -687 1222 -657 1262
rect 657 1222 687 1262
rect -781 1138 -741 1168
rect -781 168 -741 198
rect 741 1138 781 1168
rect 741 168 781 198
<< mvpsubdiffcont >>
rect -801 -1138 -761 -198
rect 761 -1138 801 -198
rect -657 -1282 657 -1242
<< mvnsubdiffcont >>
rect -657 1222 657 1262
rect -781 198 -741 1138
rect 741 198 781 1138
<< poly >>
rect -629 1168 -29 1194
rect 29 1168 629 1194
rect -629 142 -29 168
rect 29 142 629 168
rect -607 94 -51 142
rect -607 34 -587 94
rect -71 34 -51 94
rect -607 -142 -51 34
rect 51 -34 607 142
rect 51 -94 71 -34
rect 587 -94 607 -34
rect 51 -142 607 -94
rect -629 -168 -29 -142
rect 29 -168 629 -142
rect -629 -1194 -29 -1168
rect 29 -1194 629 -1168
<< polycont >>
rect -587 34 -71 94
rect 71 -94 587 -34
<< locali >>
rect -687 1222 -657 1262
rect 657 1222 687 1262
rect -781 1138 -741 1168
rect -781 168 -741 198
rect -675 1156 -641 1172
rect -675 164 -641 180
rect -17 1156 17 1172
rect -17 164 17 180
rect 641 1156 675 1172
rect 641 164 675 180
rect 741 1138 781 1168
rect 741 168 781 198
rect -607 94 -51 114
rect -607 34 -587 94
rect -71 34 -51 94
rect -607 14 -51 34
rect 51 -34 607 -14
rect 51 -94 71 -34
rect 587 -94 607 -34
rect 51 -114 607 -94
rect -801 -198 -761 -168
rect -801 -1168 -761 -1138
rect -675 -180 -641 -164
rect -675 -1172 -641 -1156
rect -17 -180 17 -164
rect -17 -1172 17 -1156
rect 641 -180 675 -164
rect 641 -1172 675 -1156
rect 761 -198 801 -168
rect 761 -1168 801 -1138
rect -687 -1282 -657 -1242
rect 657 -1282 687 -1242
<< viali >>
rect -657 1222 657 1262
rect -781 198 -741 1138
rect -675 180 -641 1156
rect -17 180 17 1156
rect 641 180 675 1156
rect 741 198 781 1138
rect -587 34 -71 94
rect 71 -94 587 -34
rect -801 -1138 -761 -198
rect -675 -1156 -641 -180
rect -17 -1156 17 -180
rect 641 -1156 675 -180
rect 761 -1138 801 -198
rect -657 -1282 657 -1242
<< metal1 >>
rect -801 1262 801 1282
rect -801 1222 -657 1262
rect 657 1222 801 1262
rect -801 1202 801 1222
rect -801 1168 -681 1202
rect 681 1168 801 1202
rect -801 1156 -635 1168
rect -801 1138 -675 1156
rect -801 198 -781 1138
rect -741 198 -675 1138
rect -801 180 -675 198
rect -641 180 -635 1156
rect -801 168 -635 180
rect -23 1156 23 1168
rect -23 180 -17 1156
rect 17 180 23 1156
rect -23 114 23 180
rect 635 1156 801 1168
rect 635 180 641 1156
rect 675 1138 801 1156
rect 675 198 741 1138
rect 781 198 801 1138
rect 675 180 801 198
rect 635 168 801 180
rect -607 94 -51 114
rect -607 34 -587 94
rect -71 34 -51 94
rect -607 14 -51 34
rect -23 14 681 114
rect 51 -34 607 -14
rect 51 -94 71 -34
rect 587 -94 607 -34
rect 51 -114 607 -94
rect -821 -180 -635 -168
rect -821 -198 -675 -180
rect -821 -1138 -801 -198
rect -761 -1138 -675 -198
rect -821 -1156 -675 -1138
rect -641 -1156 -635 -180
rect -821 -1168 -635 -1156
rect -23 -180 23 -168
rect -23 -1156 -17 -180
rect 17 -1156 23 -180
rect -23 -1168 23 -1156
rect 635 -180 681 14
rect 635 -1156 641 -180
rect 675 -1156 681 -180
rect 635 -1168 681 -1156
rect 741 -198 821 -168
rect 741 -1138 761 -198
rect 801 -1138 821 -198
rect -821 -1222 -681 -1168
rect 741 -1222 821 -1138
rect -821 -1242 821 -1222
rect -821 -1282 -657 -1242
rect 657 -1282 821 -1242
rect -821 -1302 821 -1282
<< labels >>
rlabel metal1 581 14 681 114 3 NAND
rlabel metal1 -801 1182 -701 1282 1 VDD
rlabel metal1 51 -114 607 -14 3 A
rlabel metal1 -607 14 -51 114 7 B
rlabel metal1 -821 -1302 -721 -1202 5 VSS
<< end >>
