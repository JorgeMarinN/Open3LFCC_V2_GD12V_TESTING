magic
tech sky130A
timestamp 1698272975
<< nwell >>
rect 0 0 1517 1150
<< mvpmos >>
rect 62 33 112 1117
rect 141 33 191 1117
rect 220 33 270 1117
rect 299 33 349 1117
rect 378 33 428 1117
rect 457 33 507 1117
rect 536 33 586 1117
rect 615 33 665 1117
rect 694 33 744 1117
rect 773 33 823 1117
rect 852 33 902 1117
rect 931 33 981 1117
rect 1010 33 1060 1117
rect 1089 33 1139 1117
rect 1168 33 1218 1117
rect 1247 33 1297 1117
rect 1326 33 1376 1117
rect 1405 33 1455 1117
<< mvpdiff >>
rect 33 1111 62 1117
rect 33 39 39 1111
rect 56 39 62 1111
rect 33 33 62 39
rect 112 1111 141 1117
rect 112 39 118 1111
rect 135 39 141 1111
rect 112 33 141 39
rect 191 1111 220 1117
rect 191 39 197 1111
rect 214 39 220 1111
rect 191 33 220 39
rect 270 1111 299 1117
rect 270 39 276 1111
rect 293 39 299 1111
rect 270 33 299 39
rect 349 1111 378 1117
rect 349 39 355 1111
rect 372 39 378 1111
rect 349 33 378 39
rect 428 1111 457 1117
rect 428 39 434 1111
rect 451 39 457 1111
rect 428 33 457 39
rect 507 1111 536 1117
rect 507 39 513 1111
rect 530 39 536 1111
rect 507 33 536 39
rect 586 1111 615 1117
rect 586 39 592 1111
rect 609 39 615 1111
rect 586 33 615 39
rect 665 1111 694 1117
rect 665 39 671 1111
rect 688 39 694 1111
rect 665 33 694 39
rect 744 1111 773 1117
rect 744 39 750 1111
rect 767 39 773 1111
rect 744 33 773 39
rect 823 1111 852 1117
rect 823 39 829 1111
rect 846 39 852 1111
rect 823 33 852 39
rect 902 1111 931 1117
rect 902 39 908 1111
rect 925 39 931 1111
rect 902 33 931 39
rect 981 1111 1010 1117
rect 981 39 987 1111
rect 1004 39 1010 1111
rect 981 33 1010 39
rect 1060 1111 1089 1117
rect 1060 39 1066 1111
rect 1083 39 1089 1111
rect 1060 33 1089 39
rect 1139 1111 1168 1117
rect 1139 39 1145 1111
rect 1162 39 1168 1111
rect 1139 33 1168 39
rect 1218 1111 1247 1117
rect 1218 39 1224 1111
rect 1241 39 1247 1111
rect 1218 33 1247 39
rect 1297 1111 1326 1117
rect 1297 39 1303 1111
rect 1320 39 1326 1111
rect 1297 33 1326 39
rect 1376 1111 1405 1117
rect 1376 39 1382 1111
rect 1399 39 1405 1111
rect 1376 33 1405 39
rect 1455 1111 1484 1117
rect 1455 39 1461 1111
rect 1478 39 1484 1111
rect 1455 33 1484 39
<< mvpdiffc >>
rect 39 39 56 1111
rect 118 39 135 1111
rect 197 39 214 1111
rect 276 39 293 1111
rect 355 39 372 1111
rect 434 39 451 1111
rect 513 39 530 1111
rect 592 39 609 1111
rect 671 39 688 1111
rect 750 39 767 1111
rect 829 39 846 1111
rect 908 39 925 1111
rect 987 39 1004 1111
rect 1066 39 1083 1111
rect 1145 39 1162 1111
rect 1224 39 1241 1111
rect 1303 39 1320 1111
rect 1382 39 1399 1111
rect 1461 39 1478 1111
<< poly >>
rect 62 1117 112 1130
rect 141 1117 191 1130
rect 220 1117 270 1130
rect 299 1117 349 1130
rect 378 1117 428 1130
rect 457 1117 507 1130
rect 536 1117 586 1130
rect 615 1117 665 1130
rect 694 1117 744 1130
rect 773 1117 823 1130
rect 852 1117 902 1130
rect 931 1117 981 1130
rect 1010 1117 1060 1130
rect 1089 1117 1139 1130
rect 1168 1117 1218 1130
rect 1247 1117 1297 1130
rect 1326 1117 1376 1130
rect 1405 1117 1455 1130
rect 62 20 112 33
rect 141 20 191 33
rect 220 20 270 33
rect 299 20 349 33
rect 378 20 428 33
rect 457 20 507 33
rect 536 20 586 33
rect 615 20 665 33
rect 694 20 744 33
rect 773 20 823 33
rect 852 20 902 33
rect 931 20 981 33
rect 1010 20 1060 33
rect 1089 20 1139 33
rect 1168 20 1218 33
rect 1247 20 1297 33
rect 1326 20 1376 33
rect 1405 20 1455 33
<< locali >>
rect 39 1111 56 1119
rect 39 31 56 39
rect 118 1111 135 1119
rect 118 31 135 39
rect 197 1111 214 1119
rect 197 31 214 39
rect 276 1111 293 1119
rect 276 31 293 39
rect 355 1111 372 1119
rect 355 31 372 39
rect 434 1111 451 1119
rect 434 31 451 39
rect 513 1111 530 1119
rect 513 31 530 39
rect 592 1111 609 1119
rect 592 31 609 39
rect 671 1111 688 1119
rect 671 31 688 39
rect 750 1111 767 1119
rect 750 31 767 39
rect 829 1111 846 1119
rect 829 31 846 39
rect 908 1111 925 1119
rect 908 31 925 39
rect 987 1111 1004 1119
rect 987 31 1004 39
rect 1066 1111 1083 1119
rect 1066 31 1083 39
rect 1145 1111 1162 1119
rect 1145 31 1162 39
rect 1224 1111 1241 1119
rect 1224 31 1241 39
rect 1303 1111 1320 1119
rect 1303 31 1320 39
rect 1382 1111 1399 1119
rect 1382 31 1399 39
rect 1461 1111 1478 1119
rect 1461 31 1478 39
<< viali >>
rect 39 39 56 1111
rect 118 39 135 1111
rect 197 39 214 1111
rect 276 39 293 1111
rect 355 39 372 1111
rect 434 39 451 1111
rect 513 39 530 1111
rect 592 39 609 1111
rect 671 39 688 1111
rect 750 39 767 1111
rect 829 39 846 1111
rect 908 39 925 1111
rect 987 39 1004 1111
rect 1066 39 1083 1111
rect 1145 39 1162 1111
rect 1224 39 1241 1111
rect 1303 39 1320 1111
rect 1382 39 1399 1111
rect 1461 39 1478 1111
<< metal1 >>
rect 36 1111 59 1117
rect 36 39 39 1111
rect 56 39 59 1111
rect 36 33 59 39
rect 115 1111 138 1117
rect 115 39 118 1111
rect 135 39 138 1111
rect 115 33 138 39
rect 194 1111 217 1117
rect 194 39 197 1111
rect 214 39 217 1111
rect 194 33 217 39
rect 273 1111 296 1117
rect 273 39 276 1111
rect 293 39 296 1111
rect 273 33 296 39
rect 352 1111 375 1117
rect 352 39 355 1111
rect 372 39 375 1111
rect 352 33 375 39
rect 431 1111 454 1117
rect 431 39 434 1111
rect 451 39 454 1111
rect 431 33 454 39
rect 510 1111 533 1117
rect 510 39 513 1111
rect 530 39 533 1111
rect 510 33 533 39
rect 589 1111 612 1117
rect 589 39 592 1111
rect 609 39 612 1111
rect 589 33 612 39
rect 668 1111 691 1117
rect 668 39 671 1111
rect 688 39 691 1111
rect 668 33 691 39
rect 747 1111 770 1117
rect 747 39 750 1111
rect 767 39 770 1111
rect 747 33 770 39
rect 826 1111 849 1117
rect 826 39 829 1111
rect 846 39 849 1111
rect 826 33 849 39
rect 905 1111 928 1117
rect 905 39 908 1111
rect 925 39 928 1111
rect 905 33 928 39
rect 984 1111 1007 1117
rect 984 39 987 1111
rect 1004 39 1007 1111
rect 984 33 1007 39
rect 1063 1111 1086 1117
rect 1063 39 1066 1111
rect 1083 39 1086 1111
rect 1063 33 1086 39
rect 1142 1111 1165 1117
rect 1142 39 1145 1111
rect 1162 39 1165 1111
rect 1142 33 1165 39
rect 1221 1111 1244 1117
rect 1221 39 1224 1111
rect 1241 39 1244 1111
rect 1221 33 1244 39
rect 1300 1111 1323 1117
rect 1300 39 1303 1111
rect 1320 39 1323 1111
rect 1300 33 1323 39
rect 1379 1111 1402 1117
rect 1379 39 1382 1111
rect 1399 39 1402 1111
rect 1379 33 1402 39
rect 1458 1111 1481 1117
rect 1458 39 1461 1111
rect 1478 39 1481 1111
rect 1458 33 1481 39
<< end >>
