magic
tech sky130A
timestamp 1698626380
<< mvnmos >>
rect -88 -48 -38 52
rect -9 -48 41 52
rect 70 -48 120 52
rect 149 -48 199 52
rect 228 -48 278 52
rect 307 -48 357 52
rect 386 -48 436 52
rect 465 -48 515 52
rect 544 -48 594 52
rect 623 -48 673 52
rect 702 -48 752 52
rect 781 -48 831 52
<< mvndiff >>
rect -117 46 -88 52
rect -117 -42 -111 46
rect -94 -42 -88 46
rect -117 -48 -88 -42
rect -38 46 -9 52
rect -38 -42 -32 46
rect -15 -42 -9 46
rect -38 -48 -9 -42
rect 41 46 70 52
rect 41 -42 47 46
rect 64 -42 70 46
rect 41 -48 70 -42
rect 120 46 149 52
rect 120 -42 126 46
rect 143 -42 149 46
rect 120 -48 149 -42
rect 199 46 228 52
rect 199 -42 205 46
rect 222 -42 228 46
rect 199 -48 228 -42
rect 278 46 307 52
rect 278 -42 284 46
rect 301 -42 307 46
rect 278 -48 307 -42
rect 357 46 386 52
rect 357 -42 363 46
rect 380 -42 386 46
rect 357 -48 386 -42
rect 436 46 465 52
rect 436 -42 442 46
rect 459 -42 465 46
rect 436 -48 465 -42
rect 515 46 544 52
rect 515 -42 521 46
rect 538 -42 544 46
rect 515 -48 544 -42
rect 594 46 623 52
rect 594 -42 600 46
rect 617 -42 623 46
rect 594 -48 623 -42
rect 673 46 702 52
rect 673 -42 679 46
rect 696 -42 702 46
rect 673 -48 702 -42
rect 752 46 781 52
rect 752 -42 758 46
rect 775 -42 781 46
rect 752 -48 781 -42
rect 831 46 860 52
rect 831 -42 837 46
rect 854 -42 860 46
rect 831 -48 860 -42
<< mvndiffc >>
rect -111 -42 -94 46
rect -32 -42 -15 46
rect 47 -42 64 46
rect 126 -42 143 46
rect 205 -42 222 46
rect 284 -42 301 46
rect 363 -42 380 46
rect 442 -42 459 46
rect 521 -42 538 46
rect 600 -42 617 46
rect 679 -42 696 46
rect 758 -42 775 46
rect 837 -42 854 46
<< poly >>
rect -88 52 -38 65
rect -9 52 41 65
rect 70 52 120 65
rect 149 52 199 65
rect 228 52 278 65
rect 307 52 357 65
rect 386 52 436 65
rect 465 52 515 65
rect 544 52 594 65
rect 623 52 673 65
rect 702 52 752 65
rect 781 52 831 65
rect -88 -61 -38 -48
rect -9 -61 41 -48
rect 70 -61 120 -48
rect 149 -61 199 -48
rect 228 -61 278 -48
rect 307 -61 357 -48
rect 386 -61 436 -48
rect 465 -61 515 -48
rect 544 -61 594 -48
rect 623 -61 673 -48
rect 702 -61 752 -48
rect 781 -61 831 -48
<< locali >>
rect -111 46 -94 54
rect -111 -50 -94 -42
rect -32 46 -15 54
rect -32 -50 -15 -42
rect 47 46 64 54
rect 47 -50 64 -42
rect 126 46 143 54
rect 126 -50 143 -42
rect 205 46 222 54
rect 205 -50 222 -42
rect 284 46 301 54
rect 284 -50 301 -42
rect 363 46 380 54
rect 363 -50 380 -42
rect 442 46 459 54
rect 442 -50 459 -42
rect 521 46 538 54
rect 521 -50 538 -42
rect 600 46 617 54
rect 600 -50 617 -42
rect 679 46 696 54
rect 679 -50 696 -42
rect 758 46 775 54
rect 758 -50 775 -42
rect 837 46 854 54
rect 837 -50 854 -42
<< viali >>
rect -111 -42 -94 46
rect -32 -42 -15 46
rect 47 -42 64 46
rect 126 -42 143 46
rect 205 -42 222 46
rect 284 -42 301 46
rect 363 -42 380 46
rect 442 -42 459 46
rect 521 -42 538 46
rect 600 -42 617 46
rect 679 -42 696 46
rect 758 -42 775 46
rect 837 -42 854 46
<< metal1 >>
rect -114 46 -91 52
rect -114 -42 -111 46
rect -94 -42 -91 46
rect -114 -48 -91 -42
rect -35 46 -12 52
rect -35 -42 -32 46
rect -15 -42 -12 46
rect -35 -48 -12 -42
rect 44 46 67 52
rect 44 -42 47 46
rect 64 -42 67 46
rect 44 -48 67 -42
rect 123 46 146 52
rect 123 -42 126 46
rect 143 -42 146 46
rect 123 -48 146 -42
rect 202 46 225 52
rect 202 -42 205 46
rect 222 -42 225 46
rect 202 -48 225 -42
rect 281 46 304 52
rect 281 -42 284 46
rect 301 -42 304 46
rect 281 -48 304 -42
rect 360 46 383 52
rect 360 -42 363 46
rect 380 -42 383 46
rect 360 -48 383 -42
rect 439 46 462 52
rect 439 -42 442 46
rect 459 -42 462 46
rect 439 -48 462 -42
rect 518 46 541 52
rect 518 -42 521 46
rect 538 -42 541 46
rect 518 -48 541 -42
rect 597 46 620 52
rect 597 -42 600 46
rect 617 -42 620 46
rect 597 -48 620 -42
rect 676 46 699 52
rect 676 -42 679 46
rect 696 -42 699 46
rect 676 -48 699 -42
rect 755 46 778 52
rect 755 -42 758 46
rect 775 -42 778 46
rect 755 -48 778 -42
rect 834 46 857 52
rect 834 -42 837 46
rect 854 -42 857 46
rect 834 -48 857 -42
<< end >>
