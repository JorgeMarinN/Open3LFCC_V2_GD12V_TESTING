magic
tech sky130A
timestamp 1693601183
<< checkpaint >>
rect -6555 -6605 31905 31855
<< nwell >>
rect -1125 25300 0 26425
rect 25300 25300 26475 26425
rect -1125 -1175 0 0
rect 25300 -1175 26475 0
<< pwell >>
rect -5925 26425 31275 31225
rect -5925 -1175 -1125 26425
rect 26475 -1175 31275 26425
rect -5925 -5975 31275 -1175
<< mvpmos >>
rect 25300 25331 25350 25769
rect -469 -50 -31 0
rect 25381 -50 25819 0
rect 25300 -519 25350 -81
<< mvpdiff >>
rect 25379 25769 25821 25771
rect -29 25763 0 25769
rect -29 25364 -23 25763
rect -64 25337 -23 25364
rect -6 25337 0 25763
rect -64 25331 0 25337
rect 25297 25331 25300 25769
rect 25350 25763 25821 25769
rect 25350 25337 25356 25763
rect 25373 25715 25821 25763
rect 25373 25385 25435 25715
rect 25765 25385 25821 25715
rect 25373 25337 25821 25385
rect 25350 25331 25821 25337
rect -64 25329 -31 25331
rect -469 25323 -31 25329
rect -469 25306 -463 25323
rect -37 25306 -31 25323
rect -469 25300 -31 25306
rect 25379 25329 25821 25331
rect 25381 25323 25819 25329
rect 25381 25306 25387 25323
rect 25813 25306 25819 25323
rect 25381 25300 25819 25306
rect -469 0 -31 3
rect 25381 0 25819 3
rect -469 -56 -31 -50
rect -469 -73 -463 -56
rect -37 -73 -31 -56
rect -469 -79 -31 -73
rect -471 -81 -29 -79
rect 25381 -56 25819 -50
rect 25381 -73 25387 -56
rect 25813 -73 25819 -56
rect 25381 -79 25819 -73
rect 25381 -81 25414 -79
rect -471 -87 0 -81
rect -471 -135 -23 -87
rect -471 -465 -415 -135
rect -85 -465 -23 -135
rect -471 -513 -23 -465
rect -6 -513 0 -87
rect -471 -519 0 -513
rect 25297 -519 25300 -81
rect 25350 -87 25414 -81
rect 25350 -513 25356 -87
rect 25373 -114 25414 -87
rect 25373 -513 25379 -114
rect 25350 -519 25379 -513
rect -471 -521 -29 -519
<< mvpdiffc >>
rect -23 25337 -6 25763
rect 25356 25337 25373 25763
rect -463 25306 -37 25323
rect 25387 25306 25813 25323
rect -463 -73 -37 -56
rect 25387 -73 25813 -56
rect -23 -513 -6 -87
rect 25356 -513 25373 -87
<< mvpsubdiff >>
rect -5525 30813 30875 30825
rect -5525 -5563 -5513 30813
rect -1537 26825 26887 26837
rect -1537 -1575 -1525 26825
rect 26875 -1575 26887 26825
rect -1537 -1587 26887 -1575
rect 30863 -5563 30875 30813
rect -5525 -5575 30875 -5563
<< mvnsubdiff >>
rect -1025 26313 0 26325
rect -1025 25317 -1013 26313
rect -17 26037 0 26313
rect -737 26025 0 26037
rect 25300 26313 26375 26325
rect 25300 26025 26087 26037
rect -737 25317 -725 26025
rect -1025 25300 -725 25317
rect 25435 25703 25765 25715
rect 25435 25397 25447 25703
rect 25753 25397 25765 25703
rect 25435 25385 25765 25397
rect 26075 25317 26087 26025
rect 26363 25317 26375 26313
rect 26075 25300 26375 25317
rect -1025 -1063 -1013 0
rect -737 -775 -725 0
rect -415 -147 -85 -135
rect -415 -453 -403 -147
rect -97 -453 -85 -147
rect -415 -465 -85 -453
rect 26075 -775 26087 0
rect -737 -787 0 -775
rect -17 -1063 0 -787
rect -1025 -1075 0 -1063
rect 25300 -787 26087 -775
rect 26363 -1063 26375 0
rect 25300 -1075 26375 -1063
<< mvpsubdiffcont >>
rect -5513 26837 30863 30813
rect -5513 -1587 -1537 26837
rect 26887 -1587 30863 26837
rect -5513 -5563 30863 -1587
<< mvnsubdiffcont >>
rect -1013 26037 -17 26313
rect -1013 25317 -737 26037
rect 25300 26037 26363 26313
rect 25447 25397 25753 25703
rect 26087 25317 26363 26037
rect -1013 -787 -737 0
rect -403 -453 -97 -147
rect -1013 -1063 -17 -787
rect 26087 -787 26363 0
rect 25300 -1063 26363 -787
<< poly >>
rect -550 25842 0 25850
rect -550 25808 -542 25842
rect -508 25808 0 25842
rect -550 25800 0 25808
rect 25300 25842 25900 25850
rect 25300 25808 25308 25842
rect 25342 25808 25858 25842
rect 25892 25808 25900 25842
rect 25300 25800 25900 25808
rect -550 25300 -500 25800
rect 25300 25769 25350 25800
rect 25300 25300 25350 25331
rect 25850 25300 25900 25800
rect -550 -8 -469 0
rect -550 -42 -542 -8
rect -508 -42 -469 -8
rect -550 -50 -469 -42
rect -31 -50 0 0
rect 25300 -8 25381 0
rect 25300 -42 25308 -8
rect 25342 -42 25381 -8
rect 25300 -50 25381 -42
rect 25819 -8 25900 0
rect 25819 -42 25858 -8
rect 25892 -42 25900 -8
rect 25819 -50 25900 -42
rect -550 -550 -500 -50
rect 25300 -81 25350 -50
rect 25300 -550 25350 -519
rect 25850 -550 25900 -50
rect -550 -558 0 -550
rect -550 -592 -542 -558
rect -508 -592 0 -558
rect -550 -600 0 -592
rect 25300 -558 25900 -550
rect 25300 -592 25308 -558
rect 25342 -592 25858 -558
rect 25892 -592 25900 -558
rect 25300 -600 25900 -592
<< polycont >>
rect -542 25808 -508 25842
rect 25308 25808 25342 25842
rect 25858 25808 25892 25842
rect -542 -42 -508 -8
rect 25308 -42 25342 -8
rect 25858 -42 25892 -8
rect -542 -592 -508 -558
rect 25308 -592 25342 -558
rect 25858 -592 25892 -558
<< locali >>
rect -5525 30813 30875 30825
rect -5525 -5563 -5513 30813
rect -1537 26825 26887 26837
rect -1537 -1575 -1525 26825
rect -1025 26313 0 26325
rect -1025 25317 -1013 26313
rect -17 26037 0 26313
rect -737 26025 0 26037
rect 25300 26313 26375 26325
rect 25300 26025 26087 26037
rect -737 25317 -725 26025
rect -550 25842 -500 25850
rect -550 25808 -542 25842
rect -508 25808 -500 25842
rect -550 25800 -500 25808
rect 25300 25842 25350 25850
rect 25300 25808 25308 25842
rect 25342 25808 25350 25842
rect 25300 25800 25350 25808
rect 25850 25842 25900 25850
rect 25850 25808 25858 25842
rect 25892 25808 25900 25842
rect 25850 25800 25900 25808
rect 25373 25771 25827 25777
rect -23 25763 -6 25771
rect -64 25337 -23 25364
rect -64 25329 -6 25337
rect 25356 25763 25827 25771
rect 25373 25715 25827 25763
rect 25373 25385 25435 25715
rect 25765 25385 25827 25715
rect 25373 25337 25827 25385
rect 25356 25329 25827 25337
rect -64 25323 -29 25329
rect 25373 25323 25827 25329
rect -1025 25300 -725 25317
rect -471 25306 -463 25323
rect -37 25306 -29 25323
rect 25379 25306 25387 25323
rect 25813 25306 25821 25323
rect 26075 25317 26087 26025
rect 26363 25317 26375 26313
rect 26075 25300 26375 25317
rect -1025 -1063 -1013 0
rect -737 -775 -725 0
rect -550 -8 -500 0
rect -550 -42 -542 -8
rect -508 -42 -500 -8
rect -550 -50 -500 -42
rect 25300 -8 25350 0
rect 25300 -42 25308 -8
rect 25342 -42 25350 -8
rect 25300 -50 25350 -42
rect 25850 -8 25900 0
rect 25850 -42 25858 -8
rect 25892 -42 25900 -8
rect 25850 -50 25900 -42
rect -471 -73 -463 -56
rect -37 -73 -29 -56
rect 25379 -73 25387 -56
rect 25813 -73 25821 -56
rect -477 -79 -23 -73
rect 25379 -79 25414 -73
rect -477 -87 -6 -79
rect -477 -135 -23 -87
rect -477 -465 -415 -135
rect -85 -465 -23 -135
rect -477 -513 -23 -465
rect -477 -521 -6 -513
rect 25356 -87 25414 -79
rect 25373 -114 25414 -87
rect 25356 -521 25373 -513
rect -477 -527 -23 -521
rect -550 -558 -500 -550
rect -550 -592 -542 -558
rect -508 -592 -500 -558
rect -550 -600 -500 -592
rect 25300 -558 25350 -550
rect 25300 -592 25308 -558
rect 25342 -592 25350 -558
rect 25300 -600 25350 -592
rect 25850 -558 25900 -550
rect 25850 -592 25858 -558
rect 25892 -592 25900 -558
rect 25850 -600 25900 -592
rect 26075 -775 26087 0
rect -737 -787 0 -775
rect -17 -1063 0 -787
rect -1025 -1075 0 -1063
rect 25300 -787 26087 -775
rect 26363 -1063 26375 0
rect 25300 -1075 26375 -1063
rect 26875 -1575 26887 26825
rect -1537 -1587 26887 -1575
rect 30863 -5563 30875 30813
rect -5525 -5575 30875 -5563
<< viali >>
rect -5513 26837 30863 30813
rect -5513 -1587 -1537 26837
rect -1013 26037 -19 26313
rect -1013 25319 -737 26037
rect 25300 26037 26363 26313
rect -542 25808 -508 25842
rect 25308 25808 25342 25842
rect 25858 25808 25892 25842
rect -23 25337 -6 25763
rect 25356 25337 25373 25763
rect 25435 25703 25765 25715
rect 25435 25397 25447 25703
rect 25447 25397 25753 25703
rect 25753 25397 25765 25703
rect 25435 25385 25765 25397
rect -463 25306 -37 25323
rect 25387 25306 25813 25323
rect 26087 25319 26363 26037
rect -1013 -787 -737 0
rect -542 -42 -508 -8
rect 25308 -42 25342 -8
rect 25858 -42 25892 -8
rect -463 -73 -37 -56
rect 25387 -73 25813 -56
rect -415 -147 -85 -135
rect -415 -453 -403 -147
rect -403 -453 -97 -147
rect -97 -453 -85 -147
rect -415 -465 -85 -453
rect -23 -513 -6 -87
rect 25356 -513 25373 -87
rect -542 -592 -508 -558
rect 25308 -592 25342 -558
rect 25858 -592 25892 -558
rect -1013 -1063 -19 -787
rect 26087 -787 26363 0
rect 25300 -1063 26363 -787
rect 26887 -1587 30863 26837
rect -5513 -5563 30863 -1587
<< metal1 >>
rect -5525 30813 30875 30825
rect -5525 -5563 -5513 30813
rect -1537 26825 26887 26837
rect -1537 -1575 -1525 26825
rect -1025 26313 0 26325
rect -1025 25319 -1013 26313
rect -19 26037 0 26313
rect -737 26025 0 26037
rect 25300 26313 26375 26325
rect 25300 26025 26087 26037
rect -737 25319 -725 26025
rect -550 25842 -500 25850
rect -550 25808 -542 25842
rect -508 25808 -500 25842
rect -550 25800 -500 25808
rect 25300 25842 25350 25850
rect 25300 25808 25308 25842
rect 25342 25808 25350 25842
rect 25300 25800 25350 25808
rect 25850 25842 25900 25850
rect 25850 25808 25858 25842
rect 25892 25808 25900 25842
rect 25850 25800 25900 25808
rect -474 25769 -26 25774
rect 25376 25769 25824 25774
rect -474 25763 -3 25769
rect -474 25715 -23 25763
rect -474 25385 -415 25715
rect -85 25385 -23 25715
rect -474 25337 -23 25385
rect -6 25337 -3 25763
rect -474 25331 -3 25337
rect 25353 25763 25824 25769
rect 25353 25337 25356 25763
rect 25373 25715 25824 25763
rect 25373 25385 25435 25715
rect 25765 25385 25824 25715
rect 25373 25337 25824 25385
rect 25353 25331 25824 25337
rect -474 25326 -26 25331
rect 25376 25326 25824 25331
rect -1025 25300 -725 25319
rect -469 25323 -31 25326
rect -469 25306 -463 25323
rect -37 25306 -31 25323
rect -469 25303 -31 25306
rect 25381 25323 25819 25326
rect 25381 25306 25387 25323
rect 25813 25306 25819 25323
rect 25381 25303 25819 25306
rect 26075 25319 26087 26025
rect 26363 25319 26375 26313
rect 26075 25300 26375 25319
rect -1025 -1063 -1013 0
rect -737 -775 -725 0
rect -550 -8 -500 0
rect -550 -42 -542 -8
rect -508 -42 -500 -8
rect -550 -50 -500 -42
rect 25300 -8 25350 0
rect 25300 -42 25308 -8
rect 25342 -42 25350 -8
rect 25300 -50 25350 -42
rect 25850 -8 25900 0
rect 25850 -42 25858 -8
rect 25892 -42 25900 -8
rect 25850 -50 25900 -42
rect -469 -56 -31 -53
rect -469 -73 -463 -56
rect -37 -73 -31 -56
rect -469 -76 -31 -73
rect 25381 -56 25819 -53
rect 25381 -73 25387 -56
rect 25813 -73 25819 -56
rect 25381 -76 25819 -73
rect -474 -81 -26 -76
rect 25376 -81 25824 -76
rect -474 -87 -3 -81
rect -474 -135 -23 -87
rect -474 -465 -415 -135
rect -85 -465 -23 -135
rect -474 -513 -23 -465
rect -6 -513 -3 -87
rect -474 -519 -3 -513
rect 25353 -87 25824 -81
rect 25353 -513 25356 -87
rect 25373 -135 25824 -87
rect 25373 -465 25435 -135
rect 25765 -465 25824 -135
rect 25373 -513 25824 -465
rect 25353 -519 25824 -513
rect -474 -524 -26 -519
rect 25376 -524 25824 -519
rect -550 -558 -500 -550
rect -550 -592 -542 -558
rect -508 -592 -500 -558
rect -550 -600 -500 -592
rect 25300 -558 25350 -550
rect 25300 -592 25308 -558
rect 25342 -592 25350 -558
rect 25300 -600 25350 -592
rect 25850 -558 25900 -550
rect 25850 -592 25858 -558
rect 25892 -592 25900 -558
rect 25850 -600 25900 -592
rect 26075 -775 26087 0
rect -737 -787 0 -775
rect -19 -1063 0 -787
rect -1025 -1075 0 -1063
rect 25300 -787 26087 -775
rect 26363 -1063 26375 0
rect 25300 -1075 26375 -1063
rect 26875 -1575 26887 26825
rect -1537 -1587 26887 -1575
rect 30863 -5563 30875 30813
rect -5525 -5575 30875 -5563
<< via1 >>
rect -5513 26837 30863 30813
rect -5513 1117 -1537 26825
rect 25388 26125 25488 26225
rect -542 25808 -508 25842
rect 25308 25808 25342 25842
rect 25858 25808 25892 25842
rect -415 25385 -85 25715
rect 25435 25385 25765 25715
rect 26175 25338 26275 25438
rect -925 -188 -825 -88
rect -542 -42 -508 -8
rect 25308 -42 25342 -8
rect 25858 -42 25892 -8
rect -415 -465 -85 -135
rect 25435 -465 25765 -135
rect -542 -592 -508 -558
rect 25308 -592 25342 -558
rect 25858 -592 25892 -558
rect -138 -975 -38 -875
rect 26887 -1587 30863 26837
rect -495 -5563 30863 -1587
<< metal2 >>
rect -5525 30813 30875 30825
rect -5525 26837 -5513 30813
rect -5525 26825 26887 26837
rect -5525 1117 -5513 26825
rect -1537 1117 -1525 26825
rect 25378 26225 25498 26235
rect 25378 26125 25388 26225
rect 25488 26125 25498 26225
rect 25378 26115 25498 26125
rect -725 25842 0 26025
rect -725 25808 -542 25842
rect -508 25808 0 25842
rect -725 25800 0 25808
rect 25300 25842 26075 26025
rect 25300 25808 25308 25842
rect 25342 25808 25858 25842
rect 25892 25808 26075 25842
rect 25300 25800 26075 25808
rect -725 25300 -500 25800
rect -425 25715 -75 25725
rect -425 25385 -415 25715
rect -85 25385 -75 25715
rect -425 25375 -75 25385
rect 25300 25300 25350 25800
rect 25425 25715 25775 25725
rect 25425 25385 25435 25715
rect 25765 25385 25775 25715
rect 25425 25375 25775 25385
rect 25850 25300 26075 25800
rect 26165 25438 26285 25448
rect 26165 25338 26175 25438
rect 26275 25338 26285 25438
rect 26165 25328 26285 25338
rect -725 -8 0 0
rect -725 -42 -542 -8
rect -508 -42 0 -8
rect -725 -50 0 -42
rect 25300 -8 26075 0
rect 25300 -42 25308 -8
rect 25342 -42 25858 -8
rect 25892 -42 26075 -8
rect 25300 -50 26075 -42
rect -935 -88 -815 -78
rect -935 -188 -925 -88
rect -825 -188 -815 -88
rect -935 -198 -815 -188
rect -725 -550 -500 -50
rect -425 -135 -75 -125
rect -425 -465 -415 -135
rect -85 -465 -75 -135
rect -425 -475 -75 -465
rect 25300 -550 25350 -50
rect 25425 -135 25775 -125
rect 25425 -465 25435 -135
rect 25765 -465 25775 -135
rect 25425 -475 25775 -465
rect 25850 -550 26075 -50
rect -725 -558 0 -550
rect -725 -592 -542 -558
rect -508 -592 0 -558
rect -725 -775 0 -592
rect 25300 -558 26075 -550
rect 25300 -592 25308 -558
rect 25342 -592 25858 -558
rect 25892 -592 26075 -558
rect 25300 -775 26075 -592
rect -148 -875 -28 -865
rect -148 -975 -138 -875
rect -38 -975 -28 -875
rect -148 -985 -28 -975
rect 26875 -1575 26887 26825
rect -507 -1587 26887 -1575
rect -507 -5563 -495 -1587
rect 30863 -5563 30875 30813
rect -507 -5575 30875 -5563
<< via2 >>
rect 25388 26125 25488 26225
rect -310 25490 -190 25610
rect 25540 25490 25660 25610
rect 26175 25338 26275 25438
rect -925 -188 -825 -88
rect -310 -360 -190 -240
rect 25540 -360 25660 -240
rect -138 -975 -38 -875
<< metal3 >>
rect -2525 26825 25875 27825
rect -2525 25938 -1525 26825
rect -638 25938 -186 26825
rect -2525 25614 -186 25938
rect -88 25712 0 26325
tri -186 25614 -88 25712 sw
tri -88 25624 0 25712 ne
rect 25300 26225 25664 26325
rect 25300 26125 25388 26225
rect 25488 26125 25664 26225
rect 25300 25624 25664 26125
rect -2525 25610 -88 25614
rect -2525 25490 -310 25610
rect -190 25526 -88 25610
tri -88 25526 0 25614 sw
rect -190 25490 0 25526
rect -2525 25486 0 25490
rect -2525 -575 -1525 25486
tri -412 25388 -314 25486 ne
rect -314 25388 0 25486
rect -1025 25300 -412 25388
tri -412 25300 -324 25388 sw
tri -314 25300 -226 25388 ne
rect -226 25300 0 25388
tri 25300 25526 25398 25624 ne
rect 25398 25614 25664 25624
tri 25664 25614 25762 25712 sw
rect 26875 25614 27875 25825
rect 25398 25610 27875 25614
rect 25398 25526 25540 25610
tri 25300 25438 25388 25526 sw
tri 25398 25438 25486 25526 ne
rect 25486 25490 25540 25526
rect 25660 25490 27875 25610
rect 25486 25438 27875 25490
rect 25300 25358 25388 25438
tri 25388 25358 25468 25438 sw
tri 25486 25358 25566 25438 ne
rect 25566 25358 26175 25438
rect 25300 25300 25468 25358
tri 25468 25300 25526 25358 sw
tri 25566 25300 25624 25358 ne
rect 25624 25338 26175 25358
rect 26275 25338 27875 25438
rect 25624 25300 27875 25338
rect 26875 0 27875 25300
rect -1025 -40 -324 0
tri -324 -40 -284 0 sw
tri -226 -40 -186 0 ne
rect -186 -40 0 0
rect -1025 -88 -284 -40
rect -1025 -188 -925 -88
rect -825 -138 -284 -88
tri -284 -138 -186 -40 sw
tri -186 -138 -88 -40 ne
rect -88 -138 0 -40
rect -825 -188 -186 -138
rect -1025 -236 -186 -188
tri -186 -236 -88 -138 sw
tri -88 -226 0 -138 ne
rect 25300 -40 25526 0
tri 25526 -40 25566 0 sw
tri 25624 -40 25664 0 ne
rect 25664 -40 27875 0
rect 25300 -138 25566 -40
tri 25566 -138 25664 -40 sw
tri 25664 -138 25762 -40 ne
rect 25762 -138 27875 -40
rect 25300 -226 25664 -138
rect -1025 -240 -88 -236
rect -1025 -360 -310 -240
rect -190 -324 -88 -240
tri -88 -324 0 -236 sw
rect -190 -360 0 -324
rect -1025 -364 0 -360
tri -412 -462 -314 -364 ne
rect -314 -875 0 -364
rect -314 -975 -138 -875
rect -38 -975 0 -875
rect -314 -1575 0 -975
tri 25300 -324 25398 -226 ne
rect 25398 -236 25664 -226
tri 25664 -236 25762 -138 sw
rect 25398 -240 26375 -236
rect 25398 -324 25540 -240
tri 25300 -364 25340 -324 sw
tri 25398 -364 25438 -324 ne
rect 25438 -360 25540 -324
rect 25660 -360 26375 -240
rect 25438 -364 26375 -360
rect 25300 -462 25340 -364
tri 25340 -462 25438 -364 sw
tri 25438 -462 25536 -364 ne
rect 25300 -1575 25438 -462
rect 25536 -688 26375 -364
rect 25536 -1075 25988 -688
rect 26875 -1575 27875 -138
rect -525 -2575 27875 -1575
<< via3 >>
rect 25388 26125 25488 26225
rect -310 25490 -190 25610
rect 25540 25490 25660 25610
rect 26175 25338 26275 25438
rect -925 -188 -825 -88
rect -310 -360 -190 -240
rect -138 -975 -38 -875
rect 25540 -360 25660 -240
<< metal4 >>
rect -2525 26825 25875 27825
rect -2525 25938 -1525 26825
rect -638 25938 -186 26825
rect -2525 25614 -186 25938
rect -88 25712 0 26325
tri -186 25614 -88 25712 sw
tri -88 25624 0 25712 ne
rect 25300 26225 25664 26325
rect 25300 26125 25388 26225
rect 25488 26125 25664 26225
rect 25300 25624 25664 26125
rect -2525 25610 -88 25614
rect -2525 25490 -310 25610
rect -190 25526 -88 25610
tri -88 25526 0 25614 sw
rect -190 25490 0 25526
rect -2525 25486 0 25490
rect -2525 -575 -1525 25486
tri -412 25388 -314 25486 ne
rect -314 25388 0 25486
rect -1025 25300 -412 25388
tri -412 25300 -324 25388 sw
tri -314 25300 -226 25388 ne
rect -226 25300 0 25388
tri 25300 25526 25398 25624 ne
rect 25398 25614 25664 25624
tri 25664 25614 25762 25712 sw
rect 26875 25614 27875 25825
rect 25398 25610 27875 25614
rect 25398 25526 25540 25610
tri 25300 25438 25388 25526 sw
tri 25398 25438 25486 25526 ne
rect 25486 25490 25540 25526
rect 25660 25490 27875 25610
rect 25486 25438 27875 25490
rect 25300 25358 25388 25438
tri 25388 25358 25468 25438 sw
tri 25486 25358 25566 25438 ne
rect 25566 25358 26175 25438
rect 25300 25300 25468 25358
tri 25468 25300 25526 25358 sw
tri 25566 25300 25624 25358 ne
rect 25624 25338 26175 25358
rect 26275 25338 27875 25438
rect 25624 25300 27875 25338
rect 26875 0 27875 25300
rect -1025 -40 -324 0
tri -324 -40 -284 0 sw
tri -226 -40 -186 0 ne
rect -186 -40 0 0
rect -1025 -88 -284 -40
rect -1025 -188 -925 -88
rect -825 -138 -284 -88
tri -284 -138 -186 -40 sw
tri -186 -138 -88 -40 ne
rect -88 -138 0 -40
rect -825 -188 -186 -138
rect -1025 -236 -186 -188
tri -186 -236 -88 -138 sw
tri -88 -226 0 -138 ne
rect 25300 -40 25526 0
tri 25526 -40 25566 0 sw
tri 25624 -40 25664 0 ne
rect 25664 -40 27875 0
rect 25300 -138 25566 -40
tri 25566 -138 25664 -40 sw
tri 25664 -138 25762 -40 ne
rect 25762 -138 27875 -40
rect 25300 -226 25664 -138
rect -1025 -240 -88 -236
rect -1025 -360 -310 -240
rect -190 -324 -88 -240
tri -88 -324 0 -236 sw
rect -190 -360 0 -324
rect -1025 -364 0 -360
tri -412 -462 -314 -364 ne
rect -314 -875 0 -364
rect -314 -975 -138 -875
rect -38 -975 0 -875
rect -314 -1575 0 -975
tri 25300 -324 25398 -226 ne
rect 25398 -236 25664 -226
tri 25664 -236 25762 -138 sw
rect 25398 -240 26375 -236
rect 25398 -324 25540 -240
tri 25300 -364 25340 -324 sw
tri 25398 -364 25438 -324 ne
rect 25438 -360 25540 -324
rect 25660 -360 26375 -240
rect 25438 -364 26375 -360
rect 25300 -462 25340 -364
tri 25340 -462 25438 -364 sw
tri 25438 -462 25536 -364 ne
rect 25300 -1575 25438 -462
rect 25536 -688 26375 -364
rect 25536 -1075 25988 -688
rect 26875 -1575 27875 -138
rect -525 -2575 27875 -1575
<< via4 >>
rect -310 25490 -190 25610
rect 25540 25490 25660 25610
rect -310 -360 -190 -240
rect 25540 -360 25660 -240
<< metal5 >>
rect -2525 26825 25875 27825
rect -2525 25903 -1525 26825
rect -603 25903 -292 26825
rect -2525 25610 -292 25903
tri -292 25610 -154 25748 sw
rect -53 25747 0 26325
tri -53 25694 0 25747 ne
rect 25300 25694 25558 26325
rect -2525 25592 -310 25610
rect -2525 -575 -1525 25592
tri -448 25456 -312 25592 ne
rect -312 25490 -310 25592
rect -190 25490 -154 25610
rect -312 25456 -154 25490
tri -154 25456 0 25610 sw
rect -1025 25300 -447 25353
tri -447 25300 -394 25353 sw
tri -312 25300 -156 25456 ne
rect -156 25300 0 25456
tri 25300 25456 25538 25694 ne
rect 25538 25610 25558 25694
tri 25558 25610 25696 25748 sw
rect 25538 25490 25540 25610
rect 25660 25508 25696 25610
tri 25696 25508 25798 25610 sw
rect 26875 25508 27875 25825
rect 25660 25490 27875 25508
rect 25538 25456 27875 25490
tri 25300 25300 25456 25456 sw
tri 25538 25300 25694 25456 ne
rect 25694 25300 27875 25456
rect 26875 0 27875 25300
rect -1025 -103 -394 0
tri -394 -103 -291 0 sw
tri -156 -103 -53 0 ne
rect -53 -103 0 0
rect -1025 -240 -291 -103
tri -291 -240 -154 -103 sw
tri -53 -156 0 -103 ne
rect 25300 -103 25456 0
tri 25456 -103 25559 0 sw
tri 25694 -103 25797 0 ne
rect 25797 -103 27875 0
rect 25300 -156 25559 -103
rect -1025 -258 -310 -240
tri -448 -360 -346 -258 ne
rect -346 -360 -310 -258
rect -190 -360 -154 -240
tri -346 -498 -208 -360 ne
rect -208 -394 -154 -360
tri -154 -394 0 -240 sw
rect -208 -1575 0 -394
tri 25300 -394 25538 -156 ne
rect 25538 -240 25559 -156
tri 25559 -240 25696 -103 sw
rect 25538 -360 25540 -240
rect 25660 -342 25696 -240
tri 25696 -342 25798 -240 sw
rect 25660 -360 26375 -342
rect 25538 -394 26375 -360
tri 25300 -497 25403 -394 sw
rect 25300 -1575 25403 -497
tri 25538 -498 25642 -394 ne
rect 25642 -653 26375 -394
rect 25642 -1075 25953 -653
rect 26875 -1575 27875 -103
rect -525 -2575 27875 -1575
use pmos_drain_frame_lt  pmos_drain_frame_lt_0 waffle_cells
timestamp 1675433017
transform 1 0 -550 0 1 0
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_1
timestamp 1675433017
transform 0 -1 1100 -1 0 25850
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_2
timestamp 1675433017
transform 1 0 -550 0 1 1100
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_3
timestamp 1675433017
transform 0 -1 2200 -1 0 25850
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_4
timestamp 1675433017
transform 1 0 -550 0 1 2200
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_5
timestamp 1675433017
transform 0 -1 3300 -1 0 25850
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_6
timestamp 1675433017
transform 1 0 -550 0 1 3300
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_7
timestamp 1675433017
transform 0 -1 4400 -1 0 25850
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_8
timestamp 1675433017
transform 1 0 -550 0 1 4400
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_9
timestamp 1675433017
transform 0 -1 5500 -1 0 25850
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_10
timestamp 1675433017
transform 1 0 -550 0 1 5500
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_11
timestamp 1675433017
transform 0 -1 6600 -1 0 25850
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_12
timestamp 1675433017
transform 1 0 -550 0 1 6600
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_13
timestamp 1675433017
transform 0 -1 7700 -1 0 25850
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_14
timestamp 1675433017
transform 1 0 -550 0 1 7700
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_15
timestamp 1675433017
transform 0 -1 8800 -1 0 25850
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_16
timestamp 1675433017
transform 1 0 -550 0 1 8800
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_17
timestamp 1675433017
transform 0 -1 9900 -1 0 25850
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_18
timestamp 1675433017
transform 1 0 -550 0 1 9900
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_19
timestamp 1675433017
transform 0 -1 11000 -1 0 25850
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_20
timestamp 1675433017
transform 1 0 -550 0 1 11000
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_21
timestamp 1675433017
transform 0 -1 12100 -1 0 25850
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_22
timestamp 1675433017
transform 1 0 -550 0 1 12100
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_23
timestamp 1675433017
transform 0 -1 13200 -1 0 25850
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_24
timestamp 1675433017
transform 1 0 -550 0 1 13200
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_25
timestamp 1675433017
transform 0 -1 14300 -1 0 25850
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_26
timestamp 1675433017
transform 1 0 -550 0 1 14300
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_27
timestamp 1675433017
transform 0 -1 15400 -1 0 25850
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_28
timestamp 1675433017
transform 1 0 -550 0 1 15400
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_29
timestamp 1675433017
transform 0 -1 16500 -1 0 25850
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_30
timestamp 1675433017
transform 1 0 -550 0 1 16500
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_31
timestamp 1675433017
transform 0 -1 17600 -1 0 25850
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_32
timestamp 1675433017
transform 1 0 -550 0 1 17600
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_33
timestamp 1675433017
transform 0 -1 18700 -1 0 25850
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_34
timestamp 1675433017
transform 1 0 -550 0 1 18700
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_35
timestamp 1675433017
transform 0 -1 19800 -1 0 25850
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_36
timestamp 1675433017
transform 1 0 -550 0 1 19800
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_37
timestamp 1675433017
transform 0 -1 20900 -1 0 25850
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_38
timestamp 1675433017
transform 1 0 -550 0 1 20900
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_39
timestamp 1675433017
transform 0 -1 22000 -1 0 25850
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_40
timestamp 1675433017
transform 1 0 -550 0 1 22000
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_41
timestamp 1675433017
transform 0 -1 23100 -1 0 25850
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_42
timestamp 1675433017
transform 1 0 -550 0 1 23100
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_43
timestamp 1675433017
transform 0 -1 24200 -1 0 25850
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_44
timestamp 1675433017
transform 1 0 -550 0 1 24200
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_45
timestamp 1675433017
transform 0 -1 25300 -1 0 25850
box -975 -113 663 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_0 waffle_cells
timestamp 1675433101
transform 0 -1 550 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_1
timestamp 1675433101
transform 1 0 25300 0 1 550
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_2
timestamp 1675433101
transform 0 -1 1650 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_3
timestamp 1675433101
transform 1 0 25300 0 1 1650
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_4
timestamp 1675433101
transform 0 -1 2750 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_5
timestamp 1675433101
transform 1 0 25300 0 1 2750
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_6
timestamp 1675433101
transform 0 -1 3850 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_7
timestamp 1675433101
transform 1 0 25300 0 1 3850
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_8
timestamp 1675433101
transform 0 -1 4950 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_9
timestamp 1675433101
transform 1 0 25300 0 1 4950
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_10
timestamp 1675433101
transform 0 -1 6050 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_11
timestamp 1675433101
transform 1 0 25300 0 1 6050
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_12
timestamp 1675433101
transform 0 -1 7150 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_13
timestamp 1675433101
transform 1 0 25300 0 1 7150
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_14
timestamp 1675433101
transform 0 -1 8250 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_15
timestamp 1675433101
transform 1 0 25300 0 1 8250
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_16
timestamp 1675433101
transform 0 -1 9350 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_17
timestamp 1675433101
transform 1 0 25300 0 1 9350
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_18
timestamp 1675433101
transform 0 -1 10450 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_19
timestamp 1675433101
transform 1 0 25300 0 1 10450
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_20
timestamp 1675433101
transform 0 -1 11550 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_21
timestamp 1675433101
transform 1 0 25300 0 1 11550
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_22
timestamp 1675433101
transform 0 -1 12650 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_23
timestamp 1675433101
transform 1 0 25300 0 1 12650
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_24
timestamp 1675433101
transform 0 -1 13750 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_25
timestamp 1675433101
transform 1 0 25300 0 1 13750
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_26
timestamp 1675433101
transform 0 -1 14850 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_27
timestamp 1675433101
transform 1 0 25300 0 1 14850
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_28
timestamp 1675433101
transform 0 -1 15950 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_29
timestamp 1675433101
transform 1 0 25300 0 1 15950
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_30
timestamp 1675433101
transform 0 -1 17050 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_31
timestamp 1675433101
transform 1 0 25300 0 1 17050
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_32
timestamp 1675433101
transform 0 -1 18150 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_33
timestamp 1675433101
transform 1 0 25300 0 1 18150
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_34
timestamp 1675433101
transform 0 -1 19250 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_35
timestamp 1675433101
transform 1 0 25300 0 1 19250
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_36
timestamp 1675433101
transform 0 -1 20350 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_37
timestamp 1675433101
transform 1 0 25300 0 1 20350
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_38
timestamp 1675433101
transform 0 -1 21450 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_39
timestamp 1675433101
transform 1 0 25300 0 1 21450
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_40
timestamp 1675433101
transform 0 -1 22550 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_41
timestamp 1675433101
transform 1 0 25300 0 1 22550
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_42
timestamp 1675433101
transform 0 -1 23650 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_43
timestamp 1675433101
transform 1 0 25300 0 1 23650
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_44
timestamp 1675433101
transform 0 -1 24750 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_45
timestamp 1675433101
transform 1 0 25300 0 1 24750
box -113 -113 1575 663
use pmos_drain_in  pmos_drain_in_0 waffle_cells
timestamp 1675432984
transform 1 0 0 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1
timestamp 1675432984
transform 1 0 0 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_2
timestamp 1675432984
transform 1 0 0 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_3
timestamp 1675432984
transform 1 0 0 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_4
timestamp 1675432984
transform 1 0 0 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_5
timestamp 1675432984
transform 1 0 0 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_6
timestamp 1675432984
transform 1 0 0 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_7
timestamp 1675432984
transform 1 0 0 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_8
timestamp 1675432984
transform 1 0 0 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_9
timestamp 1675432984
transform 1 0 0 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_10
timestamp 1675432984
transform 1 0 0 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_11
timestamp 1675432984
transform 1 0 0 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_12
timestamp 1675432984
transform 1 0 0 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_13
timestamp 1675432984
transform 1 0 0 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_14
timestamp 1675432984
transform 1 0 0 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_15
timestamp 1675432984
transform 1 0 0 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_16
timestamp 1675432984
transform 1 0 0 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_17
timestamp 1675432984
transform 1 0 0 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_18
timestamp 1675432984
transform 1 0 0 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_19
timestamp 1675432984
transform 1 0 0 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_20
timestamp 1675432984
transform 1 0 0 0 1 22550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_21
timestamp 1675432984
transform 1 0 0 0 1 23650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_22
timestamp 1675432984
transform 1 0 0 0 1 24750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_23
timestamp 1675432984
transform 1 0 550 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_24
timestamp 1675432984
transform 1 0 550 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_25
timestamp 1675432984
transform 1 0 550 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_26
timestamp 1675432984
transform 1 0 550 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_27
timestamp 1675432984
transform 1 0 550 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_28
timestamp 1675432984
transform 1 0 550 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_29
timestamp 1675432984
transform 1 0 550 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_30
timestamp 1675432984
transform 1 0 550 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_31
timestamp 1675432984
transform 1 0 550 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_32
timestamp 1675432984
transform 1 0 550 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_33
timestamp 1675432984
transform 1 0 550 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_34
timestamp 1675432984
transform 1 0 550 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_35
timestamp 1675432984
transform 1 0 550 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_36
timestamp 1675432984
transform 1 0 550 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_37
timestamp 1675432984
transform 1 0 550 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_38
timestamp 1675432984
transform 1 0 550 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_39
timestamp 1675432984
transform 1 0 550 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_40
timestamp 1675432984
transform 1 0 550 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_41
timestamp 1675432984
transform 1 0 550 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_42
timestamp 1675432984
transform 1 0 550 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_43
timestamp 1675432984
transform 1 0 550 0 1 22000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_44
timestamp 1675432984
transform 1 0 550 0 1 23100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_45
timestamp 1675432984
transform 1 0 550 0 1 24200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_46
timestamp 1675432984
transform 1 0 1100 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_47
timestamp 1675432984
transform 1 0 1100 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_48
timestamp 1675432984
transform 1 0 1100 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_49
timestamp 1675432984
transform 1 0 1100 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_50
timestamp 1675432984
transform 1 0 1100 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_51
timestamp 1675432984
transform 1 0 1100 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_52
timestamp 1675432984
transform 1 0 1100 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_53
timestamp 1675432984
transform 1 0 1100 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_54
timestamp 1675432984
transform 1 0 1100 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_55
timestamp 1675432984
transform 1 0 1100 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_56
timestamp 1675432984
transform 1 0 1100 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_57
timestamp 1675432984
transform 1 0 1100 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_58
timestamp 1675432984
transform 1 0 1100 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_59
timestamp 1675432984
transform 1 0 1100 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_60
timestamp 1675432984
transform 1 0 1100 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_61
timestamp 1675432984
transform 1 0 1100 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_62
timestamp 1675432984
transform 1 0 1100 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_63
timestamp 1675432984
transform 1 0 1100 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_64
timestamp 1675432984
transform 1 0 1100 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_65
timestamp 1675432984
transform 1 0 1100 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_66
timestamp 1675432984
transform 1 0 1100 0 1 22550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_67
timestamp 1675432984
transform 1 0 1100 0 1 23650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_68
timestamp 1675432984
transform 1 0 1100 0 1 24750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_69
timestamp 1675432984
transform 1 0 1650 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_70
timestamp 1675432984
transform 1 0 1650 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_71
timestamp 1675432984
transform 1 0 1650 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_72
timestamp 1675432984
transform 1 0 1650 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_73
timestamp 1675432984
transform 1 0 1650 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_74
timestamp 1675432984
transform 1 0 1650 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_75
timestamp 1675432984
transform 1 0 1650 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_76
timestamp 1675432984
transform 1 0 1650 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_77
timestamp 1675432984
transform 1 0 1650 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_78
timestamp 1675432984
transform 1 0 1650 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_79
timestamp 1675432984
transform 1 0 1650 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_80
timestamp 1675432984
transform 1 0 1650 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_81
timestamp 1675432984
transform 1 0 1650 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_82
timestamp 1675432984
transform 1 0 1650 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_83
timestamp 1675432984
transform 1 0 1650 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_84
timestamp 1675432984
transform 1 0 1650 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_85
timestamp 1675432984
transform 1 0 1650 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_86
timestamp 1675432984
transform 1 0 1650 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_87
timestamp 1675432984
transform 1 0 1650 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_88
timestamp 1675432984
transform 1 0 1650 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_89
timestamp 1675432984
transform 1 0 1650 0 1 22000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_90
timestamp 1675432984
transform 1 0 1650 0 1 23100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_91
timestamp 1675432984
transform 1 0 1650 0 1 24200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_92
timestamp 1675432984
transform 1 0 2200 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_93
timestamp 1675432984
transform 1 0 2200 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_94
timestamp 1675432984
transform 1 0 2200 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_95
timestamp 1675432984
transform 1 0 2200 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_96
timestamp 1675432984
transform 1 0 2200 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_97
timestamp 1675432984
transform 1 0 2200 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_98
timestamp 1675432984
transform 1 0 2200 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_99
timestamp 1675432984
transform 1 0 2200 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_100
timestamp 1675432984
transform 1 0 2200 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_101
timestamp 1675432984
transform 1 0 2200 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_102
timestamp 1675432984
transform 1 0 2200 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_103
timestamp 1675432984
transform 1 0 2200 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_104
timestamp 1675432984
transform 1 0 2200 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_105
timestamp 1675432984
transform 1 0 2200 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_106
timestamp 1675432984
transform 1 0 2200 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_107
timestamp 1675432984
transform 1 0 2200 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_108
timestamp 1675432984
transform 1 0 2200 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_109
timestamp 1675432984
transform 1 0 2200 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_110
timestamp 1675432984
transform 1 0 2200 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_111
timestamp 1675432984
transform 1 0 2200 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_112
timestamp 1675432984
transform 1 0 2200 0 1 22550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_113
timestamp 1675432984
transform 1 0 2200 0 1 23650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_114
timestamp 1675432984
transform 1 0 2200 0 1 24750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_115
timestamp 1675432984
transform 1 0 2750 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_116
timestamp 1675432984
transform 1 0 2750 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_117
timestamp 1675432984
transform 1 0 2750 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_118
timestamp 1675432984
transform 1 0 2750 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_119
timestamp 1675432984
transform 1 0 2750 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_120
timestamp 1675432984
transform 1 0 2750 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_121
timestamp 1675432984
transform 1 0 2750 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_122
timestamp 1675432984
transform 1 0 2750 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_123
timestamp 1675432984
transform 1 0 2750 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_124
timestamp 1675432984
transform 1 0 2750 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_125
timestamp 1675432984
transform 1 0 2750 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_126
timestamp 1675432984
transform 1 0 2750 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_127
timestamp 1675432984
transform 1 0 2750 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_128
timestamp 1675432984
transform 1 0 2750 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_129
timestamp 1675432984
transform 1 0 2750 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_130
timestamp 1675432984
transform 1 0 2750 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_131
timestamp 1675432984
transform 1 0 2750 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_132
timestamp 1675432984
transform 1 0 2750 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_133
timestamp 1675432984
transform 1 0 2750 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_134
timestamp 1675432984
transform 1 0 2750 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_135
timestamp 1675432984
transform 1 0 2750 0 1 22000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_136
timestamp 1675432984
transform 1 0 2750 0 1 23100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_137
timestamp 1675432984
transform 1 0 2750 0 1 24200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_138
timestamp 1675432984
transform 1 0 3300 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_139
timestamp 1675432984
transform 1 0 3300 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_140
timestamp 1675432984
transform 1 0 3300 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_141
timestamp 1675432984
transform 1 0 3300 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_142
timestamp 1675432984
transform 1 0 3300 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_143
timestamp 1675432984
transform 1 0 3300 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_144
timestamp 1675432984
transform 1 0 3300 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_145
timestamp 1675432984
transform 1 0 3300 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_146
timestamp 1675432984
transform 1 0 3300 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_147
timestamp 1675432984
transform 1 0 3300 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_148
timestamp 1675432984
transform 1 0 3300 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_149
timestamp 1675432984
transform 1 0 3300 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_150
timestamp 1675432984
transform 1 0 3300 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_151
timestamp 1675432984
transform 1 0 3300 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_152
timestamp 1675432984
transform 1 0 3300 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_153
timestamp 1675432984
transform 1 0 3300 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_154
timestamp 1675432984
transform 1 0 3300 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_155
timestamp 1675432984
transform 1 0 3300 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_156
timestamp 1675432984
transform 1 0 3300 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_157
timestamp 1675432984
transform 1 0 3300 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_158
timestamp 1675432984
transform 1 0 3300 0 1 22550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_159
timestamp 1675432984
transform 1 0 3300 0 1 23650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_160
timestamp 1675432984
transform 1 0 3300 0 1 24750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_161
timestamp 1675432984
transform 1 0 3850 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_162
timestamp 1675432984
transform 1 0 3850 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_163
timestamp 1675432984
transform 1 0 3850 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_164
timestamp 1675432984
transform 1 0 3850 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_165
timestamp 1675432984
transform 1 0 3850 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_166
timestamp 1675432984
transform 1 0 3850 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_167
timestamp 1675432984
transform 1 0 3850 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_168
timestamp 1675432984
transform 1 0 3850 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_169
timestamp 1675432984
transform 1 0 3850 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_170
timestamp 1675432984
transform 1 0 3850 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_171
timestamp 1675432984
transform 1 0 3850 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_172
timestamp 1675432984
transform 1 0 3850 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_173
timestamp 1675432984
transform 1 0 3850 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_174
timestamp 1675432984
transform 1 0 3850 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_175
timestamp 1675432984
transform 1 0 3850 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_176
timestamp 1675432984
transform 1 0 3850 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_177
timestamp 1675432984
transform 1 0 3850 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_178
timestamp 1675432984
transform 1 0 3850 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_179
timestamp 1675432984
transform 1 0 3850 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_180
timestamp 1675432984
transform 1 0 3850 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_181
timestamp 1675432984
transform 1 0 3850 0 1 22000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_182
timestamp 1675432984
transform 1 0 3850 0 1 23100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_183
timestamp 1675432984
transform 1 0 3850 0 1 24200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_184
timestamp 1675432984
transform 1 0 4400 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_185
timestamp 1675432984
transform 1 0 4400 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_186
timestamp 1675432984
transform 1 0 4400 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_187
timestamp 1675432984
transform 1 0 4400 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_188
timestamp 1675432984
transform 1 0 4400 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_189
timestamp 1675432984
transform 1 0 4400 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_190
timestamp 1675432984
transform 1 0 4400 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_191
timestamp 1675432984
transform 1 0 4400 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_192
timestamp 1675432984
transform 1 0 4400 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_193
timestamp 1675432984
transform 1 0 4400 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_194
timestamp 1675432984
transform 1 0 4400 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_195
timestamp 1675432984
transform 1 0 4400 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_196
timestamp 1675432984
transform 1 0 4400 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_197
timestamp 1675432984
transform 1 0 4400 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_198
timestamp 1675432984
transform 1 0 4400 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_199
timestamp 1675432984
transform 1 0 4400 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_200
timestamp 1675432984
transform 1 0 4400 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_201
timestamp 1675432984
transform 1 0 4400 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_202
timestamp 1675432984
transform 1 0 4400 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_203
timestamp 1675432984
transform 1 0 4400 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_204
timestamp 1675432984
transform 1 0 4400 0 1 22550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_205
timestamp 1675432984
transform 1 0 4400 0 1 23650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_206
timestamp 1675432984
transform 1 0 4400 0 1 24750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_207
timestamp 1675432984
transform 1 0 4950 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_208
timestamp 1675432984
transform 1 0 4950 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_209
timestamp 1675432984
transform 1 0 4950 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_210
timestamp 1675432984
transform 1 0 4950 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_211
timestamp 1675432984
transform 1 0 4950 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_212
timestamp 1675432984
transform 1 0 4950 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_213
timestamp 1675432984
transform 1 0 4950 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_214
timestamp 1675432984
transform 1 0 4950 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_215
timestamp 1675432984
transform 1 0 4950 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_216
timestamp 1675432984
transform 1 0 4950 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_217
timestamp 1675432984
transform 1 0 4950 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_218
timestamp 1675432984
transform 1 0 4950 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_219
timestamp 1675432984
transform 1 0 4950 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_220
timestamp 1675432984
transform 1 0 4950 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_221
timestamp 1675432984
transform 1 0 4950 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_222
timestamp 1675432984
transform 1 0 4950 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_223
timestamp 1675432984
transform 1 0 4950 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_224
timestamp 1675432984
transform 1 0 4950 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_225
timestamp 1675432984
transform 1 0 4950 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_226
timestamp 1675432984
transform 1 0 4950 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_227
timestamp 1675432984
transform 1 0 4950 0 1 22000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_228
timestamp 1675432984
transform 1 0 4950 0 1 23100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_229
timestamp 1675432984
transform 1 0 4950 0 1 24200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_230
timestamp 1675432984
transform 1 0 5500 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_231
timestamp 1675432984
transform 1 0 5500 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_232
timestamp 1675432984
transform 1 0 5500 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_233
timestamp 1675432984
transform 1 0 5500 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_234
timestamp 1675432984
transform 1 0 5500 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_235
timestamp 1675432984
transform 1 0 5500 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_236
timestamp 1675432984
transform 1 0 5500 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_237
timestamp 1675432984
transform 1 0 5500 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_238
timestamp 1675432984
transform 1 0 5500 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_239
timestamp 1675432984
transform 1 0 5500 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_240
timestamp 1675432984
transform 1 0 5500 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_241
timestamp 1675432984
transform 1 0 5500 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_242
timestamp 1675432984
transform 1 0 5500 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_243
timestamp 1675432984
transform 1 0 5500 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_244
timestamp 1675432984
transform 1 0 5500 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_245
timestamp 1675432984
transform 1 0 5500 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_246
timestamp 1675432984
transform 1 0 5500 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_247
timestamp 1675432984
transform 1 0 5500 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_248
timestamp 1675432984
transform 1 0 5500 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_249
timestamp 1675432984
transform 1 0 5500 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_250
timestamp 1675432984
transform 1 0 5500 0 1 22550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_251
timestamp 1675432984
transform 1 0 5500 0 1 23650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_252
timestamp 1675432984
transform 1 0 5500 0 1 24750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_253
timestamp 1675432984
transform 1 0 6050 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_254
timestamp 1675432984
transform 1 0 6050 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_255
timestamp 1675432984
transform 1 0 6050 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_256
timestamp 1675432984
transform 1 0 6050 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_257
timestamp 1675432984
transform 1 0 6050 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_258
timestamp 1675432984
transform 1 0 6050 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_259
timestamp 1675432984
transform 1 0 6050 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_260
timestamp 1675432984
transform 1 0 6050 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_261
timestamp 1675432984
transform 1 0 6050 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_262
timestamp 1675432984
transform 1 0 6050 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_263
timestamp 1675432984
transform 1 0 6050 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_264
timestamp 1675432984
transform 1 0 6050 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_265
timestamp 1675432984
transform 1 0 6050 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_266
timestamp 1675432984
transform 1 0 6050 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_267
timestamp 1675432984
transform 1 0 6050 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_268
timestamp 1675432984
transform 1 0 6050 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_269
timestamp 1675432984
transform 1 0 6050 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_270
timestamp 1675432984
transform 1 0 6050 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_271
timestamp 1675432984
transform 1 0 6050 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_272
timestamp 1675432984
transform 1 0 6050 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_273
timestamp 1675432984
transform 1 0 6050 0 1 22000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_274
timestamp 1675432984
transform 1 0 6050 0 1 23100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_275
timestamp 1675432984
transform 1 0 6050 0 1 24200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_276
timestamp 1675432984
transform 1 0 6600 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_277
timestamp 1675432984
transform 1 0 6600 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_278
timestamp 1675432984
transform 1 0 6600 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_279
timestamp 1675432984
transform 1 0 6600 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_280
timestamp 1675432984
transform 1 0 6600 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_281
timestamp 1675432984
transform 1 0 6600 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_282
timestamp 1675432984
transform 1 0 6600 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_283
timestamp 1675432984
transform 1 0 6600 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_284
timestamp 1675432984
transform 1 0 6600 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_285
timestamp 1675432984
transform 1 0 6600 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_286
timestamp 1675432984
transform 1 0 6600 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_287
timestamp 1675432984
transform 1 0 6600 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_288
timestamp 1675432984
transform 1 0 6600 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_289
timestamp 1675432984
transform 1 0 6600 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_290
timestamp 1675432984
transform 1 0 6600 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_291
timestamp 1675432984
transform 1 0 6600 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_292
timestamp 1675432984
transform 1 0 6600 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_293
timestamp 1675432984
transform 1 0 6600 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_294
timestamp 1675432984
transform 1 0 6600 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_295
timestamp 1675432984
transform 1 0 6600 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_296
timestamp 1675432984
transform 1 0 6600 0 1 22550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_297
timestamp 1675432984
transform 1 0 6600 0 1 23650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_298
timestamp 1675432984
transform 1 0 6600 0 1 24750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_299
timestamp 1675432984
transform 1 0 7150 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_300
timestamp 1675432984
transform 1 0 7150 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_301
timestamp 1675432984
transform 1 0 7150 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_302
timestamp 1675432984
transform 1 0 7150 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_303
timestamp 1675432984
transform 1 0 7150 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_304
timestamp 1675432984
transform 1 0 7150 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_305
timestamp 1675432984
transform 1 0 7150 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_306
timestamp 1675432984
transform 1 0 7150 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_307
timestamp 1675432984
transform 1 0 7150 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_308
timestamp 1675432984
transform 1 0 7150 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_309
timestamp 1675432984
transform 1 0 7150 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_310
timestamp 1675432984
transform 1 0 7150 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_311
timestamp 1675432984
transform 1 0 7150 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_312
timestamp 1675432984
transform 1 0 7150 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_313
timestamp 1675432984
transform 1 0 7150 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_314
timestamp 1675432984
transform 1 0 7150 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_315
timestamp 1675432984
transform 1 0 7150 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_316
timestamp 1675432984
transform 1 0 7150 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_317
timestamp 1675432984
transform 1 0 7150 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_318
timestamp 1675432984
transform 1 0 7150 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_319
timestamp 1675432984
transform 1 0 7150 0 1 22000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_320
timestamp 1675432984
transform 1 0 7150 0 1 23100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_321
timestamp 1675432984
transform 1 0 7150 0 1 24200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_322
timestamp 1675432984
transform 1 0 7700 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_323
timestamp 1675432984
transform 1 0 7700 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_324
timestamp 1675432984
transform 1 0 7700 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_325
timestamp 1675432984
transform 1 0 7700 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_326
timestamp 1675432984
transform 1 0 7700 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_327
timestamp 1675432984
transform 1 0 7700 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_328
timestamp 1675432984
transform 1 0 7700 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_329
timestamp 1675432984
transform 1 0 7700 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_330
timestamp 1675432984
transform 1 0 7700 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_331
timestamp 1675432984
transform 1 0 7700 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_332
timestamp 1675432984
transform 1 0 7700 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_333
timestamp 1675432984
transform 1 0 7700 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_334
timestamp 1675432984
transform 1 0 7700 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_335
timestamp 1675432984
transform 1 0 7700 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_336
timestamp 1675432984
transform 1 0 7700 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_337
timestamp 1675432984
transform 1 0 7700 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_338
timestamp 1675432984
transform 1 0 7700 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_339
timestamp 1675432984
transform 1 0 7700 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_340
timestamp 1675432984
transform 1 0 7700 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_341
timestamp 1675432984
transform 1 0 7700 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_342
timestamp 1675432984
transform 1 0 7700 0 1 22550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_343
timestamp 1675432984
transform 1 0 7700 0 1 23650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_344
timestamp 1675432984
transform 1 0 7700 0 1 24750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_345
timestamp 1675432984
transform 1 0 8250 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_346
timestamp 1675432984
transform 1 0 8250 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_347
timestamp 1675432984
transform 1 0 8250 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_348
timestamp 1675432984
transform 1 0 8250 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_349
timestamp 1675432984
transform 1 0 8250 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_350
timestamp 1675432984
transform 1 0 8250 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_351
timestamp 1675432984
transform 1 0 8250 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_352
timestamp 1675432984
transform 1 0 8250 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_353
timestamp 1675432984
transform 1 0 8250 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_354
timestamp 1675432984
transform 1 0 8250 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_355
timestamp 1675432984
transform 1 0 8250 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_356
timestamp 1675432984
transform 1 0 8250 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_357
timestamp 1675432984
transform 1 0 8250 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_358
timestamp 1675432984
transform 1 0 8250 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_359
timestamp 1675432984
transform 1 0 8250 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_360
timestamp 1675432984
transform 1 0 8250 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_361
timestamp 1675432984
transform 1 0 8250 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_362
timestamp 1675432984
transform 1 0 8250 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_363
timestamp 1675432984
transform 1 0 8250 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_364
timestamp 1675432984
transform 1 0 8250 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_365
timestamp 1675432984
transform 1 0 8250 0 1 22000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_366
timestamp 1675432984
transform 1 0 8250 0 1 23100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_367
timestamp 1675432984
transform 1 0 8250 0 1 24200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_368
timestamp 1675432984
transform 1 0 8800 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_369
timestamp 1675432984
transform 1 0 8800 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_370
timestamp 1675432984
transform 1 0 8800 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_371
timestamp 1675432984
transform 1 0 8800 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_372
timestamp 1675432984
transform 1 0 8800 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_373
timestamp 1675432984
transform 1 0 8800 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_374
timestamp 1675432984
transform 1 0 8800 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_375
timestamp 1675432984
transform 1 0 8800 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_376
timestamp 1675432984
transform 1 0 8800 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_377
timestamp 1675432984
transform 1 0 8800 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_378
timestamp 1675432984
transform 1 0 8800 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_379
timestamp 1675432984
transform 1 0 8800 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_380
timestamp 1675432984
transform 1 0 8800 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_381
timestamp 1675432984
transform 1 0 8800 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_382
timestamp 1675432984
transform 1 0 8800 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_383
timestamp 1675432984
transform 1 0 8800 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_384
timestamp 1675432984
transform 1 0 8800 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_385
timestamp 1675432984
transform 1 0 8800 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_386
timestamp 1675432984
transform 1 0 8800 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_387
timestamp 1675432984
transform 1 0 8800 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_388
timestamp 1675432984
transform 1 0 8800 0 1 22550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_389
timestamp 1675432984
transform 1 0 8800 0 1 23650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_390
timestamp 1675432984
transform 1 0 8800 0 1 24750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_391
timestamp 1675432984
transform 1 0 9350 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_392
timestamp 1675432984
transform 1 0 9350 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_393
timestamp 1675432984
transform 1 0 9350 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_394
timestamp 1675432984
transform 1 0 9350 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_395
timestamp 1675432984
transform 1 0 9350 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_396
timestamp 1675432984
transform 1 0 9350 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_397
timestamp 1675432984
transform 1 0 9350 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_398
timestamp 1675432984
transform 1 0 9350 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_399
timestamp 1675432984
transform 1 0 9350 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_400
timestamp 1675432984
transform 1 0 9350 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_401
timestamp 1675432984
transform 1 0 9350 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_402
timestamp 1675432984
transform 1 0 9350 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_403
timestamp 1675432984
transform 1 0 9350 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_404
timestamp 1675432984
transform 1 0 9350 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_405
timestamp 1675432984
transform 1 0 9350 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_406
timestamp 1675432984
transform 1 0 9350 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_407
timestamp 1675432984
transform 1 0 9350 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_408
timestamp 1675432984
transform 1 0 9350 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_409
timestamp 1675432984
transform 1 0 9350 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_410
timestamp 1675432984
transform 1 0 9350 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_411
timestamp 1675432984
transform 1 0 9350 0 1 22000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_412
timestamp 1675432984
transform 1 0 9350 0 1 23100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_413
timestamp 1675432984
transform 1 0 9350 0 1 24200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_414
timestamp 1675432984
transform 1 0 9900 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_415
timestamp 1675432984
transform 1 0 9900 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_416
timestamp 1675432984
transform 1 0 9900 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_417
timestamp 1675432984
transform 1 0 9900 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_418
timestamp 1675432984
transform 1 0 9900 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_419
timestamp 1675432984
transform 1 0 9900 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_420
timestamp 1675432984
transform 1 0 9900 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_421
timestamp 1675432984
transform 1 0 9900 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_422
timestamp 1675432984
transform 1 0 9900 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_423
timestamp 1675432984
transform 1 0 9900 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_424
timestamp 1675432984
transform 1 0 9900 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_425
timestamp 1675432984
transform 1 0 9900 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_426
timestamp 1675432984
transform 1 0 9900 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_427
timestamp 1675432984
transform 1 0 9900 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_428
timestamp 1675432984
transform 1 0 9900 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_429
timestamp 1675432984
transform 1 0 9900 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_430
timestamp 1675432984
transform 1 0 9900 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_431
timestamp 1675432984
transform 1 0 9900 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_432
timestamp 1675432984
transform 1 0 9900 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_433
timestamp 1675432984
transform 1 0 9900 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_434
timestamp 1675432984
transform 1 0 9900 0 1 22550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_435
timestamp 1675432984
transform 1 0 9900 0 1 23650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_436
timestamp 1675432984
transform 1 0 9900 0 1 24750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_437
timestamp 1675432984
transform 1 0 10450 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_438
timestamp 1675432984
transform 1 0 10450 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_439
timestamp 1675432984
transform 1 0 10450 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_440
timestamp 1675432984
transform 1 0 10450 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_441
timestamp 1675432984
transform 1 0 10450 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_442
timestamp 1675432984
transform 1 0 10450 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_443
timestamp 1675432984
transform 1 0 10450 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_444
timestamp 1675432984
transform 1 0 10450 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_445
timestamp 1675432984
transform 1 0 10450 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_446
timestamp 1675432984
transform 1 0 10450 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_447
timestamp 1675432984
transform 1 0 10450 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_448
timestamp 1675432984
transform 1 0 10450 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_449
timestamp 1675432984
transform 1 0 10450 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_450
timestamp 1675432984
transform 1 0 10450 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_451
timestamp 1675432984
transform 1 0 10450 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_452
timestamp 1675432984
transform 1 0 10450 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_453
timestamp 1675432984
transform 1 0 10450 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_454
timestamp 1675432984
transform 1 0 10450 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_455
timestamp 1675432984
transform 1 0 10450 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_456
timestamp 1675432984
transform 1 0 10450 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_457
timestamp 1675432984
transform 1 0 10450 0 1 22000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_458
timestamp 1675432984
transform 1 0 10450 0 1 23100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_459
timestamp 1675432984
transform 1 0 10450 0 1 24200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_460
timestamp 1675432984
transform 1 0 11000 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_461
timestamp 1675432984
transform 1 0 11000 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_462
timestamp 1675432984
transform 1 0 11000 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_463
timestamp 1675432984
transform 1 0 11000 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_464
timestamp 1675432984
transform 1 0 11000 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_465
timestamp 1675432984
transform 1 0 11000 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_466
timestamp 1675432984
transform 1 0 11000 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_467
timestamp 1675432984
transform 1 0 11000 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_468
timestamp 1675432984
transform 1 0 11000 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_469
timestamp 1675432984
transform 1 0 11000 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_470
timestamp 1675432984
transform 1 0 11000 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_471
timestamp 1675432984
transform 1 0 11000 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_472
timestamp 1675432984
transform 1 0 11000 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_473
timestamp 1675432984
transform 1 0 11000 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_474
timestamp 1675432984
transform 1 0 11000 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_475
timestamp 1675432984
transform 1 0 11000 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_476
timestamp 1675432984
transform 1 0 11000 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_477
timestamp 1675432984
transform 1 0 11000 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_478
timestamp 1675432984
transform 1 0 11000 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_479
timestamp 1675432984
transform 1 0 11000 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_480
timestamp 1675432984
transform 1 0 11000 0 1 22550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_481
timestamp 1675432984
transform 1 0 11000 0 1 23650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_482
timestamp 1675432984
transform 1 0 11000 0 1 24750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_483
timestamp 1675432984
transform 1 0 11550 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_484
timestamp 1675432984
transform 1 0 11550 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_485
timestamp 1675432984
transform 1 0 11550 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_486
timestamp 1675432984
transform 1 0 11550 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_487
timestamp 1675432984
transform 1 0 11550 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_488
timestamp 1675432984
transform 1 0 11550 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_489
timestamp 1675432984
transform 1 0 11550 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_490
timestamp 1675432984
transform 1 0 11550 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_491
timestamp 1675432984
transform 1 0 11550 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_492
timestamp 1675432984
transform 1 0 11550 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_493
timestamp 1675432984
transform 1 0 11550 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_494
timestamp 1675432984
transform 1 0 11550 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_495
timestamp 1675432984
transform 1 0 11550 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_496
timestamp 1675432984
transform 1 0 11550 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_497
timestamp 1675432984
transform 1 0 11550 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_498
timestamp 1675432984
transform 1 0 11550 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_499
timestamp 1675432984
transform 1 0 11550 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_500
timestamp 1675432984
transform 1 0 11550 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_501
timestamp 1675432984
transform 1 0 11550 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_502
timestamp 1675432984
transform 1 0 11550 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_503
timestamp 1675432984
transform 1 0 11550 0 1 22000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_504
timestamp 1675432984
transform 1 0 11550 0 1 23100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_505
timestamp 1675432984
transform 1 0 11550 0 1 24200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_506
timestamp 1675432984
transform 1 0 12100 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_507
timestamp 1675432984
transform 1 0 12100 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_508
timestamp 1675432984
transform 1 0 12100 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_509
timestamp 1675432984
transform 1 0 12100 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_510
timestamp 1675432984
transform 1 0 12100 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_511
timestamp 1675432984
transform 1 0 12100 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_512
timestamp 1675432984
transform 1 0 12100 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_513
timestamp 1675432984
transform 1 0 12100 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_514
timestamp 1675432984
transform 1 0 12100 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_515
timestamp 1675432984
transform 1 0 12100 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_516
timestamp 1675432984
transform 1 0 12100 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_517
timestamp 1675432984
transform 1 0 12100 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_518
timestamp 1675432984
transform 1 0 12100 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_519
timestamp 1675432984
transform 1 0 12100 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_520
timestamp 1675432984
transform 1 0 12100 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_521
timestamp 1675432984
transform 1 0 12100 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_522
timestamp 1675432984
transform 1 0 12100 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_523
timestamp 1675432984
transform 1 0 12100 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_524
timestamp 1675432984
transform 1 0 12100 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_525
timestamp 1675432984
transform 1 0 12100 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_526
timestamp 1675432984
transform 1 0 12100 0 1 22550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_527
timestamp 1675432984
transform 1 0 12100 0 1 23650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_528
timestamp 1675432984
transform 1 0 12100 0 1 24750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_529
timestamp 1675432984
transform 1 0 12650 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_530
timestamp 1675432984
transform 1 0 12650 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_531
timestamp 1675432984
transform 1 0 12650 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_532
timestamp 1675432984
transform 1 0 12650 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_533
timestamp 1675432984
transform 1 0 12650 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_534
timestamp 1675432984
transform 1 0 12650 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_535
timestamp 1675432984
transform 1 0 12650 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_536
timestamp 1675432984
transform 1 0 12650 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_537
timestamp 1675432984
transform 1 0 12650 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_538
timestamp 1675432984
transform 1 0 12650 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_539
timestamp 1675432984
transform 1 0 12650 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_540
timestamp 1675432984
transform 1 0 12650 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_541
timestamp 1675432984
transform 1 0 12650 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_542
timestamp 1675432984
transform 1 0 12650 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_543
timestamp 1675432984
transform 1 0 12650 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_544
timestamp 1675432984
transform 1 0 12650 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_545
timestamp 1675432984
transform 1 0 12650 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_546
timestamp 1675432984
transform 1 0 12650 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_547
timestamp 1675432984
transform 1 0 12650 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_548
timestamp 1675432984
transform 1 0 12650 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_549
timestamp 1675432984
transform 1 0 12650 0 1 22000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_550
timestamp 1675432984
transform 1 0 12650 0 1 23100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_551
timestamp 1675432984
transform 1 0 12650 0 1 24200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_552
timestamp 1675432984
transform 1 0 13200 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_553
timestamp 1675432984
transform 1 0 13200 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_554
timestamp 1675432984
transform 1 0 13200 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_555
timestamp 1675432984
transform 1 0 13200 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_556
timestamp 1675432984
transform 1 0 13200 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_557
timestamp 1675432984
transform 1 0 13200 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_558
timestamp 1675432984
transform 1 0 13200 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_559
timestamp 1675432984
transform 1 0 13200 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_560
timestamp 1675432984
transform 1 0 13200 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_561
timestamp 1675432984
transform 1 0 13200 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_562
timestamp 1675432984
transform 1 0 13200 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_563
timestamp 1675432984
transform 1 0 13200 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_564
timestamp 1675432984
transform 1 0 13200 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_565
timestamp 1675432984
transform 1 0 13200 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_566
timestamp 1675432984
transform 1 0 13200 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_567
timestamp 1675432984
transform 1 0 13200 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_568
timestamp 1675432984
transform 1 0 13200 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_569
timestamp 1675432984
transform 1 0 13200 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_570
timestamp 1675432984
transform 1 0 13200 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_571
timestamp 1675432984
transform 1 0 13200 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_572
timestamp 1675432984
transform 1 0 13200 0 1 22550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_573
timestamp 1675432984
transform 1 0 13200 0 1 23650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_574
timestamp 1675432984
transform 1 0 13200 0 1 24750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_575
timestamp 1675432984
transform 1 0 13750 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_576
timestamp 1675432984
transform 1 0 13750 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_577
timestamp 1675432984
transform 1 0 13750 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_578
timestamp 1675432984
transform 1 0 13750 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_579
timestamp 1675432984
transform 1 0 13750 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_580
timestamp 1675432984
transform 1 0 13750 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_581
timestamp 1675432984
transform 1 0 13750 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_582
timestamp 1675432984
transform 1 0 13750 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_583
timestamp 1675432984
transform 1 0 13750 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_584
timestamp 1675432984
transform 1 0 13750 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_585
timestamp 1675432984
transform 1 0 13750 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_586
timestamp 1675432984
transform 1 0 13750 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_587
timestamp 1675432984
transform 1 0 13750 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_588
timestamp 1675432984
transform 1 0 13750 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_589
timestamp 1675432984
transform 1 0 13750 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_590
timestamp 1675432984
transform 1 0 13750 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_591
timestamp 1675432984
transform 1 0 13750 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_592
timestamp 1675432984
transform 1 0 13750 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_593
timestamp 1675432984
transform 1 0 13750 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_594
timestamp 1675432984
transform 1 0 13750 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_595
timestamp 1675432984
transform 1 0 13750 0 1 22000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_596
timestamp 1675432984
transform 1 0 13750 0 1 23100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_597
timestamp 1675432984
transform 1 0 13750 0 1 24200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_598
timestamp 1675432984
transform 1 0 14300 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_599
timestamp 1675432984
transform 1 0 14300 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_600
timestamp 1675432984
transform 1 0 14300 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_601
timestamp 1675432984
transform 1 0 14300 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_602
timestamp 1675432984
transform 1 0 14300 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_603
timestamp 1675432984
transform 1 0 14300 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_604
timestamp 1675432984
transform 1 0 14300 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_605
timestamp 1675432984
transform 1 0 14300 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_606
timestamp 1675432984
transform 1 0 14300 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_607
timestamp 1675432984
transform 1 0 14300 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_608
timestamp 1675432984
transform 1 0 14300 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_609
timestamp 1675432984
transform 1 0 14300 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_610
timestamp 1675432984
transform 1 0 14300 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_611
timestamp 1675432984
transform 1 0 14300 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_612
timestamp 1675432984
transform 1 0 14300 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_613
timestamp 1675432984
transform 1 0 14300 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_614
timestamp 1675432984
transform 1 0 14300 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_615
timestamp 1675432984
transform 1 0 14300 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_616
timestamp 1675432984
transform 1 0 14300 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_617
timestamp 1675432984
transform 1 0 14300 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_618
timestamp 1675432984
transform 1 0 14300 0 1 22550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_619
timestamp 1675432984
transform 1 0 14300 0 1 23650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_620
timestamp 1675432984
transform 1 0 14300 0 1 24750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_621
timestamp 1675432984
transform 1 0 14850 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_622
timestamp 1675432984
transform 1 0 14850 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_623
timestamp 1675432984
transform 1 0 14850 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_624
timestamp 1675432984
transform 1 0 14850 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_625
timestamp 1675432984
transform 1 0 14850 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_626
timestamp 1675432984
transform 1 0 14850 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_627
timestamp 1675432984
transform 1 0 14850 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_628
timestamp 1675432984
transform 1 0 14850 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_629
timestamp 1675432984
transform 1 0 14850 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_630
timestamp 1675432984
transform 1 0 14850 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_631
timestamp 1675432984
transform 1 0 14850 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_632
timestamp 1675432984
transform 1 0 14850 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_633
timestamp 1675432984
transform 1 0 14850 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_634
timestamp 1675432984
transform 1 0 14850 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_635
timestamp 1675432984
transform 1 0 14850 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_636
timestamp 1675432984
transform 1 0 14850 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_637
timestamp 1675432984
transform 1 0 14850 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_638
timestamp 1675432984
transform 1 0 14850 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_639
timestamp 1675432984
transform 1 0 14850 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_640
timestamp 1675432984
transform 1 0 14850 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_641
timestamp 1675432984
transform 1 0 14850 0 1 22000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_642
timestamp 1675432984
transform 1 0 14850 0 1 23100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_643
timestamp 1675432984
transform 1 0 14850 0 1 24200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_644
timestamp 1675432984
transform 1 0 15400 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_645
timestamp 1675432984
transform 1 0 15400 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_646
timestamp 1675432984
transform 1 0 15400 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_647
timestamp 1675432984
transform 1 0 15400 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_648
timestamp 1675432984
transform 1 0 15400 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_649
timestamp 1675432984
transform 1 0 15400 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_650
timestamp 1675432984
transform 1 0 15400 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_651
timestamp 1675432984
transform 1 0 15400 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_652
timestamp 1675432984
transform 1 0 15400 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_653
timestamp 1675432984
transform 1 0 15400 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_654
timestamp 1675432984
transform 1 0 15400 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_655
timestamp 1675432984
transform 1 0 15400 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_656
timestamp 1675432984
transform 1 0 15400 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_657
timestamp 1675432984
transform 1 0 15400 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_658
timestamp 1675432984
transform 1 0 15400 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_659
timestamp 1675432984
transform 1 0 15400 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_660
timestamp 1675432984
transform 1 0 15400 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_661
timestamp 1675432984
transform 1 0 15400 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_662
timestamp 1675432984
transform 1 0 15400 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_663
timestamp 1675432984
transform 1 0 15400 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_664
timestamp 1675432984
transform 1 0 15400 0 1 22550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_665
timestamp 1675432984
transform 1 0 15400 0 1 23650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_666
timestamp 1675432984
transform 1 0 15400 0 1 24750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_667
timestamp 1675432984
transform 1 0 15950 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_668
timestamp 1675432984
transform 1 0 15950 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_669
timestamp 1675432984
transform 1 0 15950 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_670
timestamp 1675432984
transform 1 0 15950 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_671
timestamp 1675432984
transform 1 0 15950 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_672
timestamp 1675432984
transform 1 0 15950 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_673
timestamp 1675432984
transform 1 0 15950 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_674
timestamp 1675432984
transform 1 0 15950 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_675
timestamp 1675432984
transform 1 0 15950 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_676
timestamp 1675432984
transform 1 0 15950 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_677
timestamp 1675432984
transform 1 0 15950 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_678
timestamp 1675432984
transform 1 0 15950 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_679
timestamp 1675432984
transform 1 0 15950 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_680
timestamp 1675432984
transform 1 0 15950 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_681
timestamp 1675432984
transform 1 0 15950 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_682
timestamp 1675432984
transform 1 0 15950 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_683
timestamp 1675432984
transform 1 0 15950 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_684
timestamp 1675432984
transform 1 0 15950 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_685
timestamp 1675432984
transform 1 0 15950 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_686
timestamp 1675432984
transform 1 0 15950 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_687
timestamp 1675432984
transform 1 0 15950 0 1 22000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_688
timestamp 1675432984
transform 1 0 15950 0 1 23100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_689
timestamp 1675432984
transform 1 0 15950 0 1 24200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_690
timestamp 1675432984
transform 1 0 16500 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_691
timestamp 1675432984
transform 1 0 16500 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_692
timestamp 1675432984
transform 1 0 16500 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_693
timestamp 1675432984
transform 1 0 16500 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_694
timestamp 1675432984
transform 1 0 16500 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_695
timestamp 1675432984
transform 1 0 16500 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_696
timestamp 1675432984
transform 1 0 16500 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_697
timestamp 1675432984
transform 1 0 16500 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_698
timestamp 1675432984
transform 1 0 16500 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_699
timestamp 1675432984
transform 1 0 16500 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_700
timestamp 1675432984
transform 1 0 16500 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_701
timestamp 1675432984
transform 1 0 16500 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_702
timestamp 1675432984
transform 1 0 16500 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_703
timestamp 1675432984
transform 1 0 16500 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_704
timestamp 1675432984
transform 1 0 16500 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_705
timestamp 1675432984
transform 1 0 16500 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_706
timestamp 1675432984
transform 1 0 16500 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_707
timestamp 1675432984
transform 1 0 16500 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_708
timestamp 1675432984
transform 1 0 16500 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_709
timestamp 1675432984
transform 1 0 16500 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_710
timestamp 1675432984
transform 1 0 16500 0 1 22550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_711
timestamp 1675432984
transform 1 0 16500 0 1 23650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_712
timestamp 1675432984
transform 1 0 16500 0 1 24750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_713
timestamp 1675432984
transform 1 0 17050 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_714
timestamp 1675432984
transform 1 0 17050 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_715
timestamp 1675432984
transform 1 0 17050 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_716
timestamp 1675432984
transform 1 0 17050 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_717
timestamp 1675432984
transform 1 0 17050 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_718
timestamp 1675432984
transform 1 0 17050 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_719
timestamp 1675432984
transform 1 0 17050 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_720
timestamp 1675432984
transform 1 0 17050 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_721
timestamp 1675432984
transform 1 0 17050 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_722
timestamp 1675432984
transform 1 0 17050 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_723
timestamp 1675432984
transform 1 0 17050 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_724
timestamp 1675432984
transform 1 0 17050 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_725
timestamp 1675432984
transform 1 0 17050 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_726
timestamp 1675432984
transform 1 0 17050 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_727
timestamp 1675432984
transform 1 0 17050 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_728
timestamp 1675432984
transform 1 0 17050 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_729
timestamp 1675432984
transform 1 0 17050 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_730
timestamp 1675432984
transform 1 0 17050 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_731
timestamp 1675432984
transform 1 0 17050 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_732
timestamp 1675432984
transform 1 0 17050 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_733
timestamp 1675432984
transform 1 0 17050 0 1 22000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_734
timestamp 1675432984
transform 1 0 17050 0 1 23100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_735
timestamp 1675432984
transform 1 0 17050 0 1 24200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_736
timestamp 1675432984
transform 1 0 17600 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_737
timestamp 1675432984
transform 1 0 17600 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_738
timestamp 1675432984
transform 1 0 17600 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_739
timestamp 1675432984
transform 1 0 17600 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_740
timestamp 1675432984
transform 1 0 17600 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_741
timestamp 1675432984
transform 1 0 17600 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_742
timestamp 1675432984
transform 1 0 17600 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_743
timestamp 1675432984
transform 1 0 17600 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_744
timestamp 1675432984
transform 1 0 17600 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_745
timestamp 1675432984
transform 1 0 17600 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_746
timestamp 1675432984
transform 1 0 17600 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_747
timestamp 1675432984
transform 1 0 17600 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_748
timestamp 1675432984
transform 1 0 17600 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_749
timestamp 1675432984
transform 1 0 17600 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_750
timestamp 1675432984
transform 1 0 17600 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_751
timestamp 1675432984
transform 1 0 17600 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_752
timestamp 1675432984
transform 1 0 17600 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_753
timestamp 1675432984
transform 1 0 17600 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_754
timestamp 1675432984
transform 1 0 17600 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_755
timestamp 1675432984
transform 1 0 17600 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_756
timestamp 1675432984
transform 1 0 17600 0 1 22550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_757
timestamp 1675432984
transform 1 0 17600 0 1 23650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_758
timestamp 1675432984
transform 1 0 17600 0 1 24750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_759
timestamp 1675432984
transform 1 0 18150 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_760
timestamp 1675432984
transform 1 0 18150 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_761
timestamp 1675432984
transform 1 0 18150 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_762
timestamp 1675432984
transform 1 0 18150 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_763
timestamp 1675432984
transform 1 0 18150 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_764
timestamp 1675432984
transform 1 0 18150 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_765
timestamp 1675432984
transform 1 0 18150 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_766
timestamp 1675432984
transform 1 0 18150 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_767
timestamp 1675432984
transform 1 0 18150 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_768
timestamp 1675432984
transform 1 0 18150 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_769
timestamp 1675432984
transform 1 0 18150 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_770
timestamp 1675432984
transform 1 0 18150 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_771
timestamp 1675432984
transform 1 0 18150 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_772
timestamp 1675432984
transform 1 0 18150 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_773
timestamp 1675432984
transform 1 0 18150 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_774
timestamp 1675432984
transform 1 0 18150 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_775
timestamp 1675432984
transform 1 0 18150 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_776
timestamp 1675432984
transform 1 0 18150 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_777
timestamp 1675432984
transform 1 0 18150 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_778
timestamp 1675432984
transform 1 0 18150 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_779
timestamp 1675432984
transform 1 0 18150 0 1 22000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_780
timestamp 1675432984
transform 1 0 18150 0 1 23100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_781
timestamp 1675432984
transform 1 0 18150 0 1 24200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_782
timestamp 1675432984
transform 1 0 18700 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_783
timestamp 1675432984
transform 1 0 18700 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_784
timestamp 1675432984
transform 1 0 18700 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_785
timestamp 1675432984
transform 1 0 18700 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_786
timestamp 1675432984
transform 1 0 18700 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_787
timestamp 1675432984
transform 1 0 18700 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_788
timestamp 1675432984
transform 1 0 18700 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_789
timestamp 1675432984
transform 1 0 18700 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_790
timestamp 1675432984
transform 1 0 18700 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_791
timestamp 1675432984
transform 1 0 18700 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_792
timestamp 1675432984
transform 1 0 18700 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_793
timestamp 1675432984
transform 1 0 18700 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_794
timestamp 1675432984
transform 1 0 18700 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_795
timestamp 1675432984
transform 1 0 18700 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_796
timestamp 1675432984
transform 1 0 18700 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_797
timestamp 1675432984
transform 1 0 18700 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_798
timestamp 1675432984
transform 1 0 18700 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_799
timestamp 1675432984
transform 1 0 18700 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_800
timestamp 1675432984
transform 1 0 18700 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_801
timestamp 1675432984
transform 1 0 18700 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_802
timestamp 1675432984
transform 1 0 18700 0 1 22550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_803
timestamp 1675432984
transform 1 0 18700 0 1 23650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_804
timestamp 1675432984
transform 1 0 18700 0 1 24750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_805
timestamp 1675432984
transform 1 0 19250 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_806
timestamp 1675432984
transform 1 0 19250 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_807
timestamp 1675432984
transform 1 0 19250 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_808
timestamp 1675432984
transform 1 0 19250 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_809
timestamp 1675432984
transform 1 0 19250 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_810
timestamp 1675432984
transform 1 0 19250 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_811
timestamp 1675432984
transform 1 0 19250 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_812
timestamp 1675432984
transform 1 0 19250 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_813
timestamp 1675432984
transform 1 0 19250 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_814
timestamp 1675432984
transform 1 0 19250 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_815
timestamp 1675432984
transform 1 0 19250 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_816
timestamp 1675432984
transform 1 0 19250 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_817
timestamp 1675432984
transform 1 0 19250 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_818
timestamp 1675432984
transform 1 0 19250 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_819
timestamp 1675432984
transform 1 0 19250 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_820
timestamp 1675432984
transform 1 0 19250 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_821
timestamp 1675432984
transform 1 0 19250 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_822
timestamp 1675432984
transform 1 0 19250 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_823
timestamp 1675432984
transform 1 0 19250 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_824
timestamp 1675432984
transform 1 0 19250 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_825
timestamp 1675432984
transform 1 0 19250 0 1 22000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_826
timestamp 1675432984
transform 1 0 19250 0 1 23100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_827
timestamp 1675432984
transform 1 0 19250 0 1 24200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_828
timestamp 1675432984
transform 1 0 19800 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_829
timestamp 1675432984
transform 1 0 19800 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_830
timestamp 1675432984
transform 1 0 19800 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_831
timestamp 1675432984
transform 1 0 19800 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_832
timestamp 1675432984
transform 1 0 19800 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_833
timestamp 1675432984
transform 1 0 19800 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_834
timestamp 1675432984
transform 1 0 19800 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_835
timestamp 1675432984
transform 1 0 19800 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_836
timestamp 1675432984
transform 1 0 19800 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_837
timestamp 1675432984
transform 1 0 19800 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_838
timestamp 1675432984
transform 1 0 19800 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_839
timestamp 1675432984
transform 1 0 19800 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_840
timestamp 1675432984
transform 1 0 19800 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_841
timestamp 1675432984
transform 1 0 19800 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_842
timestamp 1675432984
transform 1 0 19800 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_843
timestamp 1675432984
transform 1 0 19800 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_844
timestamp 1675432984
transform 1 0 19800 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_845
timestamp 1675432984
transform 1 0 19800 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_846
timestamp 1675432984
transform 1 0 19800 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_847
timestamp 1675432984
transform 1 0 19800 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_848
timestamp 1675432984
transform 1 0 19800 0 1 22550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_849
timestamp 1675432984
transform 1 0 19800 0 1 23650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_850
timestamp 1675432984
transform 1 0 19800 0 1 24750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_851
timestamp 1675432984
transform 1 0 20350 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_852
timestamp 1675432984
transform 1 0 20350 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_853
timestamp 1675432984
transform 1 0 20350 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_854
timestamp 1675432984
transform 1 0 20350 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_855
timestamp 1675432984
transform 1 0 20350 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_856
timestamp 1675432984
transform 1 0 20350 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_857
timestamp 1675432984
transform 1 0 20350 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_858
timestamp 1675432984
transform 1 0 20350 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_859
timestamp 1675432984
transform 1 0 20350 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_860
timestamp 1675432984
transform 1 0 20350 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_861
timestamp 1675432984
transform 1 0 20350 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_862
timestamp 1675432984
transform 1 0 20350 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_863
timestamp 1675432984
transform 1 0 20350 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_864
timestamp 1675432984
transform 1 0 20350 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_865
timestamp 1675432984
transform 1 0 20350 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_866
timestamp 1675432984
transform 1 0 20350 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_867
timestamp 1675432984
transform 1 0 20350 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_868
timestamp 1675432984
transform 1 0 20350 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_869
timestamp 1675432984
transform 1 0 20350 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_870
timestamp 1675432984
transform 1 0 20350 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_871
timestamp 1675432984
transform 1 0 20350 0 1 22000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_872
timestamp 1675432984
transform 1 0 20350 0 1 23100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_873
timestamp 1675432984
transform 1 0 20350 0 1 24200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_874
timestamp 1675432984
transform 1 0 20900 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_875
timestamp 1675432984
transform 1 0 20900 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_876
timestamp 1675432984
transform 1 0 20900 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_877
timestamp 1675432984
transform 1 0 20900 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_878
timestamp 1675432984
transform 1 0 20900 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_879
timestamp 1675432984
transform 1 0 20900 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_880
timestamp 1675432984
transform 1 0 20900 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_881
timestamp 1675432984
transform 1 0 20900 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_882
timestamp 1675432984
transform 1 0 20900 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_883
timestamp 1675432984
transform 1 0 20900 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_884
timestamp 1675432984
transform 1 0 20900 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_885
timestamp 1675432984
transform 1 0 20900 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_886
timestamp 1675432984
transform 1 0 20900 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_887
timestamp 1675432984
transform 1 0 20900 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_888
timestamp 1675432984
transform 1 0 20900 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_889
timestamp 1675432984
transform 1 0 20900 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_890
timestamp 1675432984
transform 1 0 20900 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_891
timestamp 1675432984
transform 1 0 20900 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_892
timestamp 1675432984
transform 1 0 20900 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_893
timestamp 1675432984
transform 1 0 20900 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_894
timestamp 1675432984
transform 1 0 20900 0 1 22550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_895
timestamp 1675432984
transform 1 0 20900 0 1 23650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_896
timestamp 1675432984
transform 1 0 20900 0 1 24750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_897
timestamp 1675432984
transform 1 0 21450 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_898
timestamp 1675432984
transform 1 0 21450 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_899
timestamp 1675432984
transform 1 0 21450 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_900
timestamp 1675432984
transform 1 0 21450 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_901
timestamp 1675432984
transform 1 0 21450 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_902
timestamp 1675432984
transform 1 0 21450 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_903
timestamp 1675432984
transform 1 0 21450 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_904
timestamp 1675432984
transform 1 0 21450 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_905
timestamp 1675432984
transform 1 0 21450 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_906
timestamp 1675432984
transform 1 0 21450 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_907
timestamp 1675432984
transform 1 0 21450 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_908
timestamp 1675432984
transform 1 0 21450 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_909
timestamp 1675432984
transform 1 0 21450 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_910
timestamp 1675432984
transform 1 0 21450 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_911
timestamp 1675432984
transform 1 0 21450 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_912
timestamp 1675432984
transform 1 0 21450 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_913
timestamp 1675432984
transform 1 0 21450 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_914
timestamp 1675432984
transform 1 0 21450 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_915
timestamp 1675432984
transform 1 0 21450 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_916
timestamp 1675432984
transform 1 0 21450 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_917
timestamp 1675432984
transform 1 0 21450 0 1 22000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_918
timestamp 1675432984
transform 1 0 21450 0 1 23100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_919
timestamp 1675432984
transform 1 0 21450 0 1 24200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_920
timestamp 1675432984
transform 1 0 22000 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_921
timestamp 1675432984
transform 1 0 22000 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_922
timestamp 1675432984
transform 1 0 22000 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_923
timestamp 1675432984
transform 1 0 22000 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_924
timestamp 1675432984
transform 1 0 22000 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_925
timestamp 1675432984
transform 1 0 22000 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_926
timestamp 1675432984
transform 1 0 22000 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_927
timestamp 1675432984
transform 1 0 22000 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_928
timestamp 1675432984
transform 1 0 22000 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_929
timestamp 1675432984
transform 1 0 22000 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_930
timestamp 1675432984
transform 1 0 22000 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_931
timestamp 1675432984
transform 1 0 22000 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_932
timestamp 1675432984
transform 1 0 22000 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_933
timestamp 1675432984
transform 1 0 22000 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_934
timestamp 1675432984
transform 1 0 22000 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_935
timestamp 1675432984
transform 1 0 22000 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_936
timestamp 1675432984
transform 1 0 22000 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_937
timestamp 1675432984
transform 1 0 22000 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_938
timestamp 1675432984
transform 1 0 22000 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_939
timestamp 1675432984
transform 1 0 22000 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_940
timestamp 1675432984
transform 1 0 22000 0 1 22550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_941
timestamp 1675432984
transform 1 0 22000 0 1 23650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_942
timestamp 1675432984
transform 1 0 22000 0 1 24750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_943
timestamp 1675432984
transform 1 0 22550 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_944
timestamp 1675432984
transform 1 0 22550 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_945
timestamp 1675432984
transform 1 0 22550 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_946
timestamp 1675432984
transform 1 0 22550 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_947
timestamp 1675432984
transform 1 0 22550 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_948
timestamp 1675432984
transform 1 0 22550 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_949
timestamp 1675432984
transform 1 0 22550 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_950
timestamp 1675432984
transform 1 0 22550 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_951
timestamp 1675432984
transform 1 0 22550 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_952
timestamp 1675432984
transform 1 0 22550 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_953
timestamp 1675432984
transform 1 0 22550 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_954
timestamp 1675432984
transform 1 0 22550 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_955
timestamp 1675432984
transform 1 0 22550 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_956
timestamp 1675432984
transform 1 0 22550 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_957
timestamp 1675432984
transform 1 0 22550 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_958
timestamp 1675432984
transform 1 0 22550 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_959
timestamp 1675432984
transform 1 0 22550 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_960
timestamp 1675432984
transform 1 0 22550 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_961
timestamp 1675432984
transform 1 0 22550 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_962
timestamp 1675432984
transform 1 0 22550 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_963
timestamp 1675432984
transform 1 0 22550 0 1 22000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_964
timestamp 1675432984
transform 1 0 22550 0 1 23100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_965
timestamp 1675432984
transform 1 0 22550 0 1 24200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_966
timestamp 1675432984
transform 1 0 23100 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_967
timestamp 1675432984
transform 1 0 23100 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_968
timestamp 1675432984
transform 1 0 23100 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_969
timestamp 1675432984
transform 1 0 23100 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_970
timestamp 1675432984
transform 1 0 23100 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_971
timestamp 1675432984
transform 1 0 23100 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_972
timestamp 1675432984
transform 1 0 23100 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_973
timestamp 1675432984
transform 1 0 23100 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_974
timestamp 1675432984
transform 1 0 23100 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_975
timestamp 1675432984
transform 1 0 23100 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_976
timestamp 1675432984
transform 1 0 23100 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_977
timestamp 1675432984
transform 1 0 23100 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_978
timestamp 1675432984
transform 1 0 23100 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_979
timestamp 1675432984
transform 1 0 23100 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_980
timestamp 1675432984
transform 1 0 23100 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_981
timestamp 1675432984
transform 1 0 23100 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_982
timestamp 1675432984
transform 1 0 23100 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_983
timestamp 1675432984
transform 1 0 23100 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_984
timestamp 1675432984
transform 1 0 23100 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_985
timestamp 1675432984
transform 1 0 23100 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_986
timestamp 1675432984
transform 1 0 23100 0 1 22550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_987
timestamp 1675432984
transform 1 0 23100 0 1 23650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_988
timestamp 1675432984
transform 1 0 23100 0 1 24750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_989
timestamp 1675432984
transform 1 0 23650 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_990
timestamp 1675432984
transform 1 0 23650 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_991
timestamp 1675432984
transform 1 0 23650 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_992
timestamp 1675432984
transform 1 0 23650 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_993
timestamp 1675432984
transform 1 0 23650 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_994
timestamp 1675432984
transform 1 0 23650 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_995
timestamp 1675432984
transform 1 0 23650 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_996
timestamp 1675432984
transform 1 0 23650 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_997
timestamp 1675432984
transform 1 0 23650 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_998
timestamp 1675432984
transform 1 0 23650 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_999
timestamp 1675432984
transform 1 0 23650 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1000
timestamp 1675432984
transform 1 0 23650 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1001
timestamp 1675432984
transform 1 0 23650 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1002
timestamp 1675432984
transform 1 0 23650 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1003
timestamp 1675432984
transform 1 0 23650 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1004
timestamp 1675432984
transform 1 0 23650 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1005
timestamp 1675432984
transform 1 0 23650 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1006
timestamp 1675432984
transform 1 0 23650 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1007
timestamp 1675432984
transform 1 0 23650 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1008
timestamp 1675432984
transform 1 0 23650 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1009
timestamp 1675432984
transform 1 0 23650 0 1 22000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1010
timestamp 1675432984
transform 1 0 23650 0 1 23100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1011
timestamp 1675432984
transform 1 0 23650 0 1 24200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1012
timestamp 1675432984
transform 1 0 24200 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1013
timestamp 1675432984
transform 1 0 24200 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1014
timestamp 1675432984
transform 1 0 24200 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1015
timestamp 1675432984
transform 1 0 24200 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1016
timestamp 1675432984
transform 1 0 24200 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1017
timestamp 1675432984
transform 1 0 24200 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1018
timestamp 1675432984
transform 1 0 24200 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1019
timestamp 1675432984
transform 1 0 24200 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1020
timestamp 1675432984
transform 1 0 24200 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1021
timestamp 1675432984
transform 1 0 24200 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1022
timestamp 1675432984
transform 1 0 24200 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1023
timestamp 1675432984
transform 1 0 24200 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1024
timestamp 1675432984
transform 1 0 24200 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1025
timestamp 1675432984
transform 1 0 24200 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1026
timestamp 1675432984
transform 1 0 24200 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1027
timestamp 1675432984
transform 1 0 24200 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1028
timestamp 1675432984
transform 1 0 24200 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1029
timestamp 1675432984
transform 1 0 24200 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1030
timestamp 1675432984
transform 1 0 24200 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1031
timestamp 1675432984
transform 1 0 24200 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1032
timestamp 1675432984
transform 1 0 24200 0 1 22550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1033
timestamp 1675432984
transform 1 0 24200 0 1 23650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1034
timestamp 1675432984
transform 1 0 24200 0 1 24750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1035
timestamp 1675432984
transform 1 0 24750 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1036
timestamp 1675432984
transform 1 0 24750 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1037
timestamp 1675432984
transform 1 0 24750 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1038
timestamp 1675432984
transform 1 0 24750 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1039
timestamp 1675432984
transform 1 0 24750 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1040
timestamp 1675432984
transform 1 0 24750 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1041
timestamp 1675432984
transform 1 0 24750 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1042
timestamp 1675432984
transform 1 0 24750 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1043
timestamp 1675432984
transform 1 0 24750 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1044
timestamp 1675432984
transform 1 0 24750 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1045
timestamp 1675432984
transform 1 0 24750 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1046
timestamp 1675432984
transform 1 0 24750 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1047
timestamp 1675432984
transform 1 0 24750 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1048
timestamp 1675432984
transform 1 0 24750 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1049
timestamp 1675432984
transform 1 0 24750 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1050
timestamp 1675432984
transform 1 0 24750 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1051
timestamp 1675432984
transform 1 0 24750 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1052
timestamp 1675432984
transform 1 0 24750 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1053
timestamp 1675432984
transform 1 0 24750 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1054
timestamp 1675432984
transform 1 0 24750 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1055
timestamp 1675432984
transform 1 0 24750 0 1 22000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1056
timestamp 1675432984
transform 1 0 24750 0 1 23100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1057
timestamp 1675432984
transform 1 0 24750 0 1 24200
box -113 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_0 waffle_cells
timestamp 1675433049
transform 0 -1 550 -1 0 25850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_1
timestamp 1675433049
transform 1 0 -550 0 1 550
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_2
timestamp 1675433049
transform 0 -1 1650 -1 0 25850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_3
timestamp 1675433049
transform 1 0 -550 0 1 1650
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_4
timestamp 1675433049
transform 0 -1 2750 -1 0 25850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_5
timestamp 1675433049
transform 1 0 -550 0 1 2750
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_6
timestamp 1675433049
transform 0 -1 3850 -1 0 25850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_7
timestamp 1675433049
transform 1 0 -550 0 1 3850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_8
timestamp 1675433049
transform 0 -1 4950 -1 0 25850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_9
timestamp 1675433049
transform 1 0 -550 0 1 4950
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_10
timestamp 1675433049
transform 0 -1 6050 -1 0 25850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_11
timestamp 1675433049
transform 1 0 -550 0 1 6050
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_12
timestamp 1675433049
transform 0 -1 7150 -1 0 25850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_13
timestamp 1675433049
transform 1 0 -550 0 1 7150
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_14
timestamp 1675433049
transform 0 -1 8250 -1 0 25850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_15
timestamp 1675433049
transform 1 0 -550 0 1 8250
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_16
timestamp 1675433049
transform 0 -1 9350 -1 0 25850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_17
timestamp 1675433049
transform 1 0 -550 0 1 9350
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_18
timestamp 1675433049
transform 0 -1 10450 -1 0 25850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_19
timestamp 1675433049
transform 1 0 -550 0 1 10450
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_20
timestamp 1675433049
transform 0 -1 11550 -1 0 25850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_21
timestamp 1675433049
transform 1 0 -550 0 1 11550
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_22
timestamp 1675433049
transform 0 -1 12650 -1 0 25850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_23
timestamp 1675433049
transform 1 0 -550 0 1 12650
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_24
timestamp 1675433049
transform 0 -1 13750 -1 0 25850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_25
timestamp 1675433049
transform 1 0 -550 0 1 13750
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_26
timestamp 1675433049
transform 0 -1 14850 -1 0 25850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_27
timestamp 1675433049
transform 1 0 -550 0 1 14850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_28
timestamp 1675433049
transform 0 -1 15950 -1 0 25850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_29
timestamp 1675433049
transform 1 0 -550 0 1 15950
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_30
timestamp 1675433049
transform 0 -1 17050 -1 0 25850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_31
timestamp 1675433049
transform 1 0 -550 0 1 17050
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_32
timestamp 1675433049
transform 0 -1 18150 -1 0 25850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_33
timestamp 1675433049
transform 1 0 -550 0 1 18150
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_34
timestamp 1675433049
transform 0 -1 19250 -1 0 25850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_35
timestamp 1675433049
transform 1 0 -550 0 1 19250
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_36
timestamp 1675433049
transform 0 -1 20350 -1 0 25850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_37
timestamp 1675433049
transform 1 0 -550 0 1 20350
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_38
timestamp 1675433049
transform 0 -1 21450 -1 0 25850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_39
timestamp 1675433049
transform 1 0 -550 0 1 21450
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_40
timestamp 1675433049
transform 0 -1 22550 -1 0 25850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_41
timestamp 1675433049
transform 1 0 -550 0 1 22550
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_42
timestamp 1675433049
transform 0 -1 23650 -1 0 25850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_43
timestamp 1675433049
transform 1 0 -550 0 1 23650
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_44
timestamp 1675433049
transform 0 -1 24750 -1 0 25850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_45
timestamp 1675433049
transform 1 0 -550 0 1 24750
box -975 -113 663 663
use pmos_source_frame_rb  pmos_source_frame_rb_0 waffle_cells
timestamp 1675433193
transform 1 0 25300 0 1 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_1
timestamp 1675433193
transform 0 -1 1100 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_2
timestamp 1675433193
transform 1 0 25300 0 1 1100
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_3
timestamp 1675433193
transform 0 -1 2200 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_4
timestamp 1675433193
transform 1 0 25300 0 1 2200
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_5
timestamp 1675433193
transform 0 -1 3300 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_6
timestamp 1675433193
transform 1 0 25300 0 1 3300
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_7
timestamp 1675433193
transform 0 -1 4400 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_8
timestamp 1675433193
transform 1 0 25300 0 1 4400
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_9
timestamp 1675433193
transform 0 -1 5500 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_10
timestamp 1675433193
transform 1 0 25300 0 1 5500
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_11
timestamp 1675433193
transform 0 -1 6600 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_12
timestamp 1675433193
transform 1 0 25300 0 1 6600
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_13
timestamp 1675433193
transform 0 -1 7700 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_14
timestamp 1675433193
transform 1 0 25300 0 1 7700
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_15
timestamp 1675433193
transform 0 -1 8800 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_16
timestamp 1675433193
transform 1 0 25300 0 1 8800
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_17
timestamp 1675433193
transform 0 -1 9900 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_18
timestamp 1675433193
transform 1 0 25300 0 1 9900
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_19
timestamp 1675433193
transform 0 -1 11000 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_20
timestamp 1675433193
transform 1 0 25300 0 1 11000
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_21
timestamp 1675433193
transform 0 -1 12100 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_22
timestamp 1675433193
transform 1 0 25300 0 1 12100
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_23
timestamp 1675433193
transform 0 -1 13200 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_24
timestamp 1675433193
transform 1 0 25300 0 1 13200
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_25
timestamp 1675433193
transform 0 -1 14300 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_26
timestamp 1675433193
transform 1 0 25300 0 1 14300
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_27
timestamp 1675433193
transform 0 -1 15400 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_28
timestamp 1675433193
transform 1 0 25300 0 1 15400
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_29
timestamp 1675433193
transform 0 -1 16500 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_30
timestamp 1675433193
transform 1 0 25300 0 1 16500
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_31
timestamp 1675433193
transform 0 -1 17600 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_32
timestamp 1675433193
transform 1 0 25300 0 1 17600
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_33
timestamp 1675433193
transform 0 -1 18700 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_34
timestamp 1675433193
transform 1 0 25300 0 1 18700
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_35
timestamp 1675433193
transform 0 -1 19800 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_36
timestamp 1675433193
transform 1 0 25300 0 1 19800
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_37
timestamp 1675433193
transform 0 -1 20900 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_38
timestamp 1675433193
transform 1 0 25300 0 1 20900
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_39
timestamp 1675433193
transform 0 -1 22000 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_40
timestamp 1675433193
transform 1 0 25300 0 1 22000
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_41
timestamp 1675433193
transform 0 -1 23100 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_42
timestamp 1675433193
transform 1 0 25300 0 1 23100
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_43
timestamp 1675433193
transform 0 -1 24200 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_44
timestamp 1675433193
transform 1 0 25300 0 1 24200
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_45
timestamp 1675433193
transform 0 -1 25300 -1 0 0
box -113 -113 1575 663
use pmos_source_in  pmos_source_in_0 waffle_cells
timestamp 1675432918
transform 1 0 0 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1
timestamp 1675432918
transform 1 0 0 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_2
timestamp 1675432918
transform 1 0 0 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_3
timestamp 1675432918
transform 1 0 0 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_4
timestamp 1675432918
transform 1 0 0 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_5
timestamp 1675432918
transform 1 0 0 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_6
timestamp 1675432918
transform 1 0 0 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_7
timestamp 1675432918
transform 1 0 0 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_8
timestamp 1675432918
transform 1 0 0 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_9
timestamp 1675432918
transform 1 0 0 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_10
timestamp 1675432918
transform 1 0 0 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_11
timestamp 1675432918
transform 1 0 0 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_12
timestamp 1675432918
transform 1 0 0 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_13
timestamp 1675432918
transform 1 0 0 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_14
timestamp 1675432918
transform 1 0 0 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_15
timestamp 1675432918
transform 1 0 0 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_16
timestamp 1675432918
transform 1 0 0 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_17
timestamp 1675432918
transform 1 0 0 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_18
timestamp 1675432918
transform 1 0 0 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_19
timestamp 1675432918
transform 1 0 0 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_20
timestamp 1675432918
transform 1 0 0 0 1 22000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_21
timestamp 1675432918
transform 1 0 0 0 1 23100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_22
timestamp 1675432918
transform 1 0 0 0 1 24200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_23
timestamp 1675432918
transform 1 0 550 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_24
timestamp 1675432918
transform 1 0 550 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_25
timestamp 1675432918
transform 1 0 550 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_26
timestamp 1675432918
transform 1 0 550 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_27
timestamp 1675432918
transform 1 0 550 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_28
timestamp 1675432918
transform 1 0 550 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_29
timestamp 1675432918
transform 1 0 550 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_30
timestamp 1675432918
transform 1 0 550 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_31
timestamp 1675432918
transform 1 0 550 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_32
timestamp 1675432918
transform 1 0 550 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_33
timestamp 1675432918
transform 1 0 550 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_34
timestamp 1675432918
transform 1 0 550 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_35
timestamp 1675432918
transform 1 0 550 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_36
timestamp 1675432918
transform 1 0 550 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_37
timestamp 1675432918
transform 1 0 550 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_38
timestamp 1675432918
transform 1 0 550 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_39
timestamp 1675432918
transform 1 0 550 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_40
timestamp 1675432918
transform 1 0 550 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_41
timestamp 1675432918
transform 1 0 550 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_42
timestamp 1675432918
transform 1 0 550 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_43
timestamp 1675432918
transform 1 0 550 0 1 22550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_44
timestamp 1675432918
transform 1 0 550 0 1 23650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_45
timestamp 1675432918
transform 1 0 550 0 1 24750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_46
timestamp 1675432918
transform 1 0 1100 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_47
timestamp 1675432918
transform 1 0 1100 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_48
timestamp 1675432918
transform 1 0 1100 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_49
timestamp 1675432918
transform 1 0 1100 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_50
timestamp 1675432918
transform 1 0 1100 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_51
timestamp 1675432918
transform 1 0 1100 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_52
timestamp 1675432918
transform 1 0 1100 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_53
timestamp 1675432918
transform 1 0 1100 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_54
timestamp 1675432918
transform 1 0 1100 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_55
timestamp 1675432918
transform 1 0 1100 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_56
timestamp 1675432918
transform 1 0 1100 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_57
timestamp 1675432918
transform 1 0 1100 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_58
timestamp 1675432918
transform 1 0 1100 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_59
timestamp 1675432918
transform 1 0 1100 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_60
timestamp 1675432918
transform 1 0 1100 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_61
timestamp 1675432918
transform 1 0 1100 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_62
timestamp 1675432918
transform 1 0 1100 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_63
timestamp 1675432918
transform 1 0 1100 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_64
timestamp 1675432918
transform 1 0 1100 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_65
timestamp 1675432918
transform 1 0 1100 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_66
timestamp 1675432918
transform 1 0 1100 0 1 22000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_67
timestamp 1675432918
transform 1 0 1100 0 1 23100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_68
timestamp 1675432918
transform 1 0 1100 0 1 24200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_69
timestamp 1675432918
transform 1 0 1650 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_70
timestamp 1675432918
transform 1 0 1650 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_71
timestamp 1675432918
transform 1 0 1650 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_72
timestamp 1675432918
transform 1 0 1650 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_73
timestamp 1675432918
transform 1 0 1650 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_74
timestamp 1675432918
transform 1 0 1650 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_75
timestamp 1675432918
transform 1 0 1650 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_76
timestamp 1675432918
transform 1 0 1650 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_77
timestamp 1675432918
transform 1 0 1650 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_78
timestamp 1675432918
transform 1 0 1650 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_79
timestamp 1675432918
transform 1 0 1650 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_80
timestamp 1675432918
transform 1 0 1650 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_81
timestamp 1675432918
transform 1 0 1650 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_82
timestamp 1675432918
transform 1 0 1650 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_83
timestamp 1675432918
transform 1 0 1650 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_84
timestamp 1675432918
transform 1 0 1650 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_85
timestamp 1675432918
transform 1 0 1650 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_86
timestamp 1675432918
transform 1 0 1650 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_87
timestamp 1675432918
transform 1 0 1650 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_88
timestamp 1675432918
transform 1 0 1650 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_89
timestamp 1675432918
transform 1 0 1650 0 1 22550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_90
timestamp 1675432918
transform 1 0 1650 0 1 23650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_91
timestamp 1675432918
transform 1 0 1650 0 1 24750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_92
timestamp 1675432918
transform 1 0 2200 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_93
timestamp 1675432918
transform 1 0 2200 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_94
timestamp 1675432918
transform 1 0 2200 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_95
timestamp 1675432918
transform 1 0 2200 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_96
timestamp 1675432918
transform 1 0 2200 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_97
timestamp 1675432918
transform 1 0 2200 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_98
timestamp 1675432918
transform 1 0 2200 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_99
timestamp 1675432918
transform 1 0 2200 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_100
timestamp 1675432918
transform 1 0 2200 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_101
timestamp 1675432918
transform 1 0 2200 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_102
timestamp 1675432918
transform 1 0 2200 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_103
timestamp 1675432918
transform 1 0 2200 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_104
timestamp 1675432918
transform 1 0 2200 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_105
timestamp 1675432918
transform 1 0 2200 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_106
timestamp 1675432918
transform 1 0 2200 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_107
timestamp 1675432918
transform 1 0 2200 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_108
timestamp 1675432918
transform 1 0 2200 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_109
timestamp 1675432918
transform 1 0 2200 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_110
timestamp 1675432918
transform 1 0 2200 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_111
timestamp 1675432918
transform 1 0 2200 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_112
timestamp 1675432918
transform 1 0 2200 0 1 22000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_113
timestamp 1675432918
transform 1 0 2200 0 1 23100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_114
timestamp 1675432918
transform 1 0 2200 0 1 24200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_115
timestamp 1675432918
transform 1 0 2750 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_116
timestamp 1675432918
transform 1 0 2750 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_117
timestamp 1675432918
transform 1 0 2750 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_118
timestamp 1675432918
transform 1 0 2750 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_119
timestamp 1675432918
transform 1 0 2750 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_120
timestamp 1675432918
transform 1 0 2750 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_121
timestamp 1675432918
transform 1 0 2750 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_122
timestamp 1675432918
transform 1 0 2750 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_123
timestamp 1675432918
transform 1 0 2750 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_124
timestamp 1675432918
transform 1 0 2750 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_125
timestamp 1675432918
transform 1 0 2750 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_126
timestamp 1675432918
transform 1 0 2750 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_127
timestamp 1675432918
transform 1 0 2750 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_128
timestamp 1675432918
transform 1 0 2750 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_129
timestamp 1675432918
transform 1 0 2750 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_130
timestamp 1675432918
transform 1 0 2750 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_131
timestamp 1675432918
transform 1 0 2750 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_132
timestamp 1675432918
transform 1 0 2750 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_133
timestamp 1675432918
transform 1 0 2750 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_134
timestamp 1675432918
transform 1 0 2750 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_135
timestamp 1675432918
transform 1 0 2750 0 1 22550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_136
timestamp 1675432918
transform 1 0 2750 0 1 23650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_137
timestamp 1675432918
transform 1 0 2750 0 1 24750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_138
timestamp 1675432918
transform 1 0 3300 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_139
timestamp 1675432918
transform 1 0 3300 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_140
timestamp 1675432918
transform 1 0 3300 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_141
timestamp 1675432918
transform 1 0 3300 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_142
timestamp 1675432918
transform 1 0 3300 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_143
timestamp 1675432918
transform 1 0 3300 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_144
timestamp 1675432918
transform 1 0 3300 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_145
timestamp 1675432918
transform 1 0 3300 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_146
timestamp 1675432918
transform 1 0 3300 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_147
timestamp 1675432918
transform 1 0 3300 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_148
timestamp 1675432918
transform 1 0 3300 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_149
timestamp 1675432918
transform 1 0 3300 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_150
timestamp 1675432918
transform 1 0 3300 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_151
timestamp 1675432918
transform 1 0 3300 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_152
timestamp 1675432918
transform 1 0 3300 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_153
timestamp 1675432918
transform 1 0 3300 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_154
timestamp 1675432918
transform 1 0 3300 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_155
timestamp 1675432918
transform 1 0 3300 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_156
timestamp 1675432918
transform 1 0 3300 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_157
timestamp 1675432918
transform 1 0 3300 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_158
timestamp 1675432918
transform 1 0 3300 0 1 22000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_159
timestamp 1675432918
transform 1 0 3300 0 1 23100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_160
timestamp 1675432918
transform 1 0 3300 0 1 24200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_161
timestamp 1675432918
transform 1 0 3850 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_162
timestamp 1675432918
transform 1 0 3850 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_163
timestamp 1675432918
transform 1 0 3850 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_164
timestamp 1675432918
transform 1 0 3850 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_165
timestamp 1675432918
transform 1 0 3850 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_166
timestamp 1675432918
transform 1 0 3850 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_167
timestamp 1675432918
transform 1 0 3850 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_168
timestamp 1675432918
transform 1 0 3850 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_169
timestamp 1675432918
transform 1 0 3850 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_170
timestamp 1675432918
transform 1 0 3850 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_171
timestamp 1675432918
transform 1 0 3850 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_172
timestamp 1675432918
transform 1 0 3850 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_173
timestamp 1675432918
transform 1 0 3850 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_174
timestamp 1675432918
transform 1 0 3850 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_175
timestamp 1675432918
transform 1 0 3850 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_176
timestamp 1675432918
transform 1 0 3850 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_177
timestamp 1675432918
transform 1 0 3850 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_178
timestamp 1675432918
transform 1 0 3850 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_179
timestamp 1675432918
transform 1 0 3850 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_180
timestamp 1675432918
transform 1 0 3850 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_181
timestamp 1675432918
transform 1 0 3850 0 1 22550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_182
timestamp 1675432918
transform 1 0 3850 0 1 23650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_183
timestamp 1675432918
transform 1 0 3850 0 1 24750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_184
timestamp 1675432918
transform 1 0 4400 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_185
timestamp 1675432918
transform 1 0 4400 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_186
timestamp 1675432918
transform 1 0 4400 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_187
timestamp 1675432918
transform 1 0 4400 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_188
timestamp 1675432918
transform 1 0 4400 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_189
timestamp 1675432918
transform 1 0 4400 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_190
timestamp 1675432918
transform 1 0 4400 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_191
timestamp 1675432918
transform 1 0 4400 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_192
timestamp 1675432918
transform 1 0 4400 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_193
timestamp 1675432918
transform 1 0 4400 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_194
timestamp 1675432918
transform 1 0 4400 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_195
timestamp 1675432918
transform 1 0 4400 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_196
timestamp 1675432918
transform 1 0 4400 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_197
timestamp 1675432918
transform 1 0 4400 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_198
timestamp 1675432918
transform 1 0 4400 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_199
timestamp 1675432918
transform 1 0 4400 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_200
timestamp 1675432918
transform 1 0 4400 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_201
timestamp 1675432918
transform 1 0 4400 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_202
timestamp 1675432918
transform 1 0 4400 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_203
timestamp 1675432918
transform 1 0 4400 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_204
timestamp 1675432918
transform 1 0 4400 0 1 22000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_205
timestamp 1675432918
transform 1 0 4400 0 1 23100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_206
timestamp 1675432918
transform 1 0 4400 0 1 24200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_207
timestamp 1675432918
transform 1 0 4950 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_208
timestamp 1675432918
transform 1 0 4950 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_209
timestamp 1675432918
transform 1 0 4950 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_210
timestamp 1675432918
transform 1 0 4950 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_211
timestamp 1675432918
transform 1 0 4950 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_212
timestamp 1675432918
transform 1 0 4950 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_213
timestamp 1675432918
transform 1 0 4950 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_214
timestamp 1675432918
transform 1 0 4950 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_215
timestamp 1675432918
transform 1 0 4950 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_216
timestamp 1675432918
transform 1 0 4950 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_217
timestamp 1675432918
transform 1 0 4950 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_218
timestamp 1675432918
transform 1 0 4950 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_219
timestamp 1675432918
transform 1 0 4950 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_220
timestamp 1675432918
transform 1 0 4950 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_221
timestamp 1675432918
transform 1 0 4950 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_222
timestamp 1675432918
transform 1 0 4950 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_223
timestamp 1675432918
transform 1 0 4950 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_224
timestamp 1675432918
transform 1 0 4950 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_225
timestamp 1675432918
transform 1 0 4950 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_226
timestamp 1675432918
transform 1 0 4950 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_227
timestamp 1675432918
transform 1 0 4950 0 1 22550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_228
timestamp 1675432918
transform 1 0 4950 0 1 23650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_229
timestamp 1675432918
transform 1 0 4950 0 1 24750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_230
timestamp 1675432918
transform 1 0 5500 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_231
timestamp 1675432918
transform 1 0 5500 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_232
timestamp 1675432918
transform 1 0 5500 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_233
timestamp 1675432918
transform 1 0 5500 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_234
timestamp 1675432918
transform 1 0 5500 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_235
timestamp 1675432918
transform 1 0 5500 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_236
timestamp 1675432918
transform 1 0 5500 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_237
timestamp 1675432918
transform 1 0 5500 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_238
timestamp 1675432918
transform 1 0 5500 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_239
timestamp 1675432918
transform 1 0 5500 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_240
timestamp 1675432918
transform 1 0 5500 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_241
timestamp 1675432918
transform 1 0 5500 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_242
timestamp 1675432918
transform 1 0 5500 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_243
timestamp 1675432918
transform 1 0 5500 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_244
timestamp 1675432918
transform 1 0 5500 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_245
timestamp 1675432918
transform 1 0 5500 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_246
timestamp 1675432918
transform 1 0 5500 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_247
timestamp 1675432918
transform 1 0 5500 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_248
timestamp 1675432918
transform 1 0 5500 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_249
timestamp 1675432918
transform 1 0 5500 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_250
timestamp 1675432918
transform 1 0 5500 0 1 22000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_251
timestamp 1675432918
transform 1 0 5500 0 1 23100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_252
timestamp 1675432918
transform 1 0 5500 0 1 24200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_253
timestamp 1675432918
transform 1 0 6050 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_254
timestamp 1675432918
transform 1 0 6050 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_255
timestamp 1675432918
transform 1 0 6050 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_256
timestamp 1675432918
transform 1 0 6050 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_257
timestamp 1675432918
transform 1 0 6050 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_258
timestamp 1675432918
transform 1 0 6050 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_259
timestamp 1675432918
transform 1 0 6050 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_260
timestamp 1675432918
transform 1 0 6050 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_261
timestamp 1675432918
transform 1 0 6050 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_262
timestamp 1675432918
transform 1 0 6050 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_263
timestamp 1675432918
transform 1 0 6050 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_264
timestamp 1675432918
transform 1 0 6050 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_265
timestamp 1675432918
transform 1 0 6050 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_266
timestamp 1675432918
transform 1 0 6050 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_267
timestamp 1675432918
transform 1 0 6050 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_268
timestamp 1675432918
transform 1 0 6050 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_269
timestamp 1675432918
transform 1 0 6050 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_270
timestamp 1675432918
transform 1 0 6050 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_271
timestamp 1675432918
transform 1 0 6050 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_272
timestamp 1675432918
transform 1 0 6050 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_273
timestamp 1675432918
transform 1 0 6050 0 1 22550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_274
timestamp 1675432918
transform 1 0 6050 0 1 23650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_275
timestamp 1675432918
transform 1 0 6050 0 1 24750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_276
timestamp 1675432918
transform 1 0 6600 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_277
timestamp 1675432918
transform 1 0 6600 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_278
timestamp 1675432918
transform 1 0 6600 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_279
timestamp 1675432918
transform 1 0 6600 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_280
timestamp 1675432918
transform 1 0 6600 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_281
timestamp 1675432918
transform 1 0 6600 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_282
timestamp 1675432918
transform 1 0 6600 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_283
timestamp 1675432918
transform 1 0 6600 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_284
timestamp 1675432918
transform 1 0 6600 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_285
timestamp 1675432918
transform 1 0 6600 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_286
timestamp 1675432918
transform 1 0 6600 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_287
timestamp 1675432918
transform 1 0 6600 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_288
timestamp 1675432918
transform 1 0 6600 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_289
timestamp 1675432918
transform 1 0 6600 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_290
timestamp 1675432918
transform 1 0 6600 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_291
timestamp 1675432918
transform 1 0 6600 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_292
timestamp 1675432918
transform 1 0 6600 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_293
timestamp 1675432918
transform 1 0 6600 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_294
timestamp 1675432918
transform 1 0 6600 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_295
timestamp 1675432918
transform 1 0 6600 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_296
timestamp 1675432918
transform 1 0 6600 0 1 22000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_297
timestamp 1675432918
transform 1 0 6600 0 1 23100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_298
timestamp 1675432918
transform 1 0 6600 0 1 24200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_299
timestamp 1675432918
transform 1 0 7150 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_300
timestamp 1675432918
transform 1 0 7150 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_301
timestamp 1675432918
transform 1 0 7150 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_302
timestamp 1675432918
transform 1 0 7150 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_303
timestamp 1675432918
transform 1 0 7150 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_304
timestamp 1675432918
transform 1 0 7150 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_305
timestamp 1675432918
transform 1 0 7150 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_306
timestamp 1675432918
transform 1 0 7150 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_307
timestamp 1675432918
transform 1 0 7150 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_308
timestamp 1675432918
transform 1 0 7150 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_309
timestamp 1675432918
transform 1 0 7150 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_310
timestamp 1675432918
transform 1 0 7150 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_311
timestamp 1675432918
transform 1 0 7150 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_312
timestamp 1675432918
transform 1 0 7150 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_313
timestamp 1675432918
transform 1 0 7150 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_314
timestamp 1675432918
transform 1 0 7150 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_315
timestamp 1675432918
transform 1 0 7150 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_316
timestamp 1675432918
transform 1 0 7150 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_317
timestamp 1675432918
transform 1 0 7150 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_318
timestamp 1675432918
transform 1 0 7150 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_319
timestamp 1675432918
transform 1 0 7150 0 1 22550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_320
timestamp 1675432918
transform 1 0 7150 0 1 23650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_321
timestamp 1675432918
transform 1 0 7150 0 1 24750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_322
timestamp 1675432918
transform 1 0 7700 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_323
timestamp 1675432918
transform 1 0 7700 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_324
timestamp 1675432918
transform 1 0 7700 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_325
timestamp 1675432918
transform 1 0 7700 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_326
timestamp 1675432918
transform 1 0 7700 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_327
timestamp 1675432918
transform 1 0 7700 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_328
timestamp 1675432918
transform 1 0 7700 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_329
timestamp 1675432918
transform 1 0 7700 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_330
timestamp 1675432918
transform 1 0 7700 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_331
timestamp 1675432918
transform 1 0 7700 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_332
timestamp 1675432918
transform 1 0 7700 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_333
timestamp 1675432918
transform 1 0 7700 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_334
timestamp 1675432918
transform 1 0 7700 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_335
timestamp 1675432918
transform 1 0 7700 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_336
timestamp 1675432918
transform 1 0 7700 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_337
timestamp 1675432918
transform 1 0 7700 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_338
timestamp 1675432918
transform 1 0 7700 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_339
timestamp 1675432918
transform 1 0 7700 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_340
timestamp 1675432918
transform 1 0 7700 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_341
timestamp 1675432918
transform 1 0 7700 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_342
timestamp 1675432918
transform 1 0 7700 0 1 22000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_343
timestamp 1675432918
transform 1 0 7700 0 1 23100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_344
timestamp 1675432918
transform 1 0 7700 0 1 24200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_345
timestamp 1675432918
transform 1 0 8250 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_346
timestamp 1675432918
transform 1 0 8250 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_347
timestamp 1675432918
transform 1 0 8250 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_348
timestamp 1675432918
transform 1 0 8250 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_349
timestamp 1675432918
transform 1 0 8250 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_350
timestamp 1675432918
transform 1 0 8250 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_351
timestamp 1675432918
transform 1 0 8250 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_352
timestamp 1675432918
transform 1 0 8250 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_353
timestamp 1675432918
transform 1 0 8250 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_354
timestamp 1675432918
transform 1 0 8250 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_355
timestamp 1675432918
transform 1 0 8250 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_356
timestamp 1675432918
transform 1 0 8250 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_357
timestamp 1675432918
transform 1 0 8250 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_358
timestamp 1675432918
transform 1 0 8250 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_359
timestamp 1675432918
transform 1 0 8250 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_360
timestamp 1675432918
transform 1 0 8250 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_361
timestamp 1675432918
transform 1 0 8250 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_362
timestamp 1675432918
transform 1 0 8250 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_363
timestamp 1675432918
transform 1 0 8250 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_364
timestamp 1675432918
transform 1 0 8250 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_365
timestamp 1675432918
transform 1 0 8250 0 1 22550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_366
timestamp 1675432918
transform 1 0 8250 0 1 23650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_367
timestamp 1675432918
transform 1 0 8250 0 1 24750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_368
timestamp 1675432918
transform 1 0 8800 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_369
timestamp 1675432918
transform 1 0 8800 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_370
timestamp 1675432918
transform 1 0 8800 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_371
timestamp 1675432918
transform 1 0 8800 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_372
timestamp 1675432918
transform 1 0 8800 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_373
timestamp 1675432918
transform 1 0 8800 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_374
timestamp 1675432918
transform 1 0 8800 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_375
timestamp 1675432918
transform 1 0 8800 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_376
timestamp 1675432918
transform 1 0 8800 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_377
timestamp 1675432918
transform 1 0 8800 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_378
timestamp 1675432918
transform 1 0 8800 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_379
timestamp 1675432918
transform 1 0 8800 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_380
timestamp 1675432918
transform 1 0 8800 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_381
timestamp 1675432918
transform 1 0 8800 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_382
timestamp 1675432918
transform 1 0 8800 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_383
timestamp 1675432918
transform 1 0 8800 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_384
timestamp 1675432918
transform 1 0 8800 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_385
timestamp 1675432918
transform 1 0 8800 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_386
timestamp 1675432918
transform 1 0 8800 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_387
timestamp 1675432918
transform 1 0 8800 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_388
timestamp 1675432918
transform 1 0 8800 0 1 22000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_389
timestamp 1675432918
transform 1 0 8800 0 1 23100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_390
timestamp 1675432918
transform 1 0 8800 0 1 24200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_391
timestamp 1675432918
transform 1 0 9350 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_392
timestamp 1675432918
transform 1 0 9350 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_393
timestamp 1675432918
transform 1 0 9350 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_394
timestamp 1675432918
transform 1 0 9350 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_395
timestamp 1675432918
transform 1 0 9350 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_396
timestamp 1675432918
transform 1 0 9350 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_397
timestamp 1675432918
transform 1 0 9350 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_398
timestamp 1675432918
transform 1 0 9350 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_399
timestamp 1675432918
transform 1 0 9350 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_400
timestamp 1675432918
transform 1 0 9350 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_401
timestamp 1675432918
transform 1 0 9350 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_402
timestamp 1675432918
transform 1 0 9350 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_403
timestamp 1675432918
transform 1 0 9350 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_404
timestamp 1675432918
transform 1 0 9350 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_405
timestamp 1675432918
transform 1 0 9350 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_406
timestamp 1675432918
transform 1 0 9350 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_407
timestamp 1675432918
transform 1 0 9350 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_408
timestamp 1675432918
transform 1 0 9350 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_409
timestamp 1675432918
transform 1 0 9350 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_410
timestamp 1675432918
transform 1 0 9350 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_411
timestamp 1675432918
transform 1 0 9350 0 1 22550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_412
timestamp 1675432918
transform 1 0 9350 0 1 23650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_413
timestamp 1675432918
transform 1 0 9350 0 1 24750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_414
timestamp 1675432918
transform 1 0 9900 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_415
timestamp 1675432918
transform 1 0 9900 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_416
timestamp 1675432918
transform 1 0 9900 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_417
timestamp 1675432918
transform 1 0 9900 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_418
timestamp 1675432918
transform 1 0 9900 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_419
timestamp 1675432918
transform 1 0 9900 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_420
timestamp 1675432918
transform 1 0 9900 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_421
timestamp 1675432918
transform 1 0 9900 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_422
timestamp 1675432918
transform 1 0 9900 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_423
timestamp 1675432918
transform 1 0 9900 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_424
timestamp 1675432918
transform 1 0 9900 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_425
timestamp 1675432918
transform 1 0 9900 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_426
timestamp 1675432918
transform 1 0 9900 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_427
timestamp 1675432918
transform 1 0 9900 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_428
timestamp 1675432918
transform 1 0 9900 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_429
timestamp 1675432918
transform 1 0 9900 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_430
timestamp 1675432918
transform 1 0 9900 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_431
timestamp 1675432918
transform 1 0 9900 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_432
timestamp 1675432918
transform 1 0 9900 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_433
timestamp 1675432918
transform 1 0 9900 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_434
timestamp 1675432918
transform 1 0 9900 0 1 22000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_435
timestamp 1675432918
transform 1 0 9900 0 1 23100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_436
timestamp 1675432918
transform 1 0 9900 0 1 24200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_437
timestamp 1675432918
transform 1 0 10450 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_438
timestamp 1675432918
transform 1 0 10450 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_439
timestamp 1675432918
transform 1 0 10450 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_440
timestamp 1675432918
transform 1 0 10450 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_441
timestamp 1675432918
transform 1 0 10450 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_442
timestamp 1675432918
transform 1 0 10450 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_443
timestamp 1675432918
transform 1 0 10450 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_444
timestamp 1675432918
transform 1 0 10450 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_445
timestamp 1675432918
transform 1 0 10450 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_446
timestamp 1675432918
transform 1 0 10450 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_447
timestamp 1675432918
transform 1 0 10450 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_448
timestamp 1675432918
transform 1 0 10450 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_449
timestamp 1675432918
transform 1 0 10450 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_450
timestamp 1675432918
transform 1 0 10450 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_451
timestamp 1675432918
transform 1 0 10450 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_452
timestamp 1675432918
transform 1 0 10450 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_453
timestamp 1675432918
transform 1 0 10450 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_454
timestamp 1675432918
transform 1 0 10450 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_455
timestamp 1675432918
transform 1 0 10450 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_456
timestamp 1675432918
transform 1 0 10450 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_457
timestamp 1675432918
transform 1 0 10450 0 1 22550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_458
timestamp 1675432918
transform 1 0 10450 0 1 23650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_459
timestamp 1675432918
transform 1 0 10450 0 1 24750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_460
timestamp 1675432918
transform 1 0 11000 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_461
timestamp 1675432918
transform 1 0 11000 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_462
timestamp 1675432918
transform 1 0 11000 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_463
timestamp 1675432918
transform 1 0 11000 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_464
timestamp 1675432918
transform 1 0 11000 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_465
timestamp 1675432918
transform 1 0 11000 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_466
timestamp 1675432918
transform 1 0 11000 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_467
timestamp 1675432918
transform 1 0 11000 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_468
timestamp 1675432918
transform 1 0 11000 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_469
timestamp 1675432918
transform 1 0 11000 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_470
timestamp 1675432918
transform 1 0 11000 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_471
timestamp 1675432918
transform 1 0 11000 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_472
timestamp 1675432918
transform 1 0 11000 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_473
timestamp 1675432918
transform 1 0 11000 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_474
timestamp 1675432918
transform 1 0 11000 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_475
timestamp 1675432918
transform 1 0 11000 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_476
timestamp 1675432918
transform 1 0 11000 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_477
timestamp 1675432918
transform 1 0 11000 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_478
timestamp 1675432918
transform 1 0 11000 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_479
timestamp 1675432918
transform 1 0 11000 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_480
timestamp 1675432918
transform 1 0 11000 0 1 22000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_481
timestamp 1675432918
transform 1 0 11000 0 1 23100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_482
timestamp 1675432918
transform 1 0 11000 0 1 24200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_483
timestamp 1675432918
transform 1 0 11550 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_484
timestamp 1675432918
transform 1 0 11550 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_485
timestamp 1675432918
transform 1 0 11550 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_486
timestamp 1675432918
transform 1 0 11550 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_487
timestamp 1675432918
transform 1 0 11550 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_488
timestamp 1675432918
transform 1 0 11550 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_489
timestamp 1675432918
transform 1 0 11550 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_490
timestamp 1675432918
transform 1 0 11550 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_491
timestamp 1675432918
transform 1 0 11550 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_492
timestamp 1675432918
transform 1 0 11550 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_493
timestamp 1675432918
transform 1 0 11550 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_494
timestamp 1675432918
transform 1 0 11550 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_495
timestamp 1675432918
transform 1 0 11550 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_496
timestamp 1675432918
transform 1 0 11550 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_497
timestamp 1675432918
transform 1 0 11550 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_498
timestamp 1675432918
transform 1 0 11550 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_499
timestamp 1675432918
transform 1 0 11550 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_500
timestamp 1675432918
transform 1 0 11550 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_501
timestamp 1675432918
transform 1 0 11550 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_502
timestamp 1675432918
transform 1 0 11550 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_503
timestamp 1675432918
transform 1 0 11550 0 1 22550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_504
timestamp 1675432918
transform 1 0 11550 0 1 23650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_505
timestamp 1675432918
transform 1 0 11550 0 1 24750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_506
timestamp 1675432918
transform 1 0 12100 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_507
timestamp 1675432918
transform 1 0 12100 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_508
timestamp 1675432918
transform 1 0 12100 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_509
timestamp 1675432918
transform 1 0 12100 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_510
timestamp 1675432918
transform 1 0 12100 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_511
timestamp 1675432918
transform 1 0 12100 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_512
timestamp 1675432918
transform 1 0 12100 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_513
timestamp 1675432918
transform 1 0 12100 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_514
timestamp 1675432918
transform 1 0 12100 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_515
timestamp 1675432918
transform 1 0 12100 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_516
timestamp 1675432918
transform 1 0 12100 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_517
timestamp 1675432918
transform 1 0 12100 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_518
timestamp 1675432918
transform 1 0 12100 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_519
timestamp 1675432918
transform 1 0 12100 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_520
timestamp 1675432918
transform 1 0 12100 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_521
timestamp 1675432918
transform 1 0 12100 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_522
timestamp 1675432918
transform 1 0 12100 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_523
timestamp 1675432918
transform 1 0 12100 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_524
timestamp 1675432918
transform 1 0 12100 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_525
timestamp 1675432918
transform 1 0 12100 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_526
timestamp 1675432918
transform 1 0 12100 0 1 22000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_527
timestamp 1675432918
transform 1 0 12100 0 1 23100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_528
timestamp 1675432918
transform 1 0 12100 0 1 24200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_529
timestamp 1675432918
transform 1 0 12650 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_530
timestamp 1675432918
transform 1 0 12650 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_531
timestamp 1675432918
transform 1 0 12650 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_532
timestamp 1675432918
transform 1 0 12650 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_533
timestamp 1675432918
transform 1 0 12650 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_534
timestamp 1675432918
transform 1 0 12650 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_535
timestamp 1675432918
transform 1 0 12650 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_536
timestamp 1675432918
transform 1 0 12650 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_537
timestamp 1675432918
transform 1 0 12650 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_538
timestamp 1675432918
transform 1 0 12650 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_539
timestamp 1675432918
transform 1 0 12650 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_540
timestamp 1675432918
transform 1 0 12650 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_541
timestamp 1675432918
transform 1 0 12650 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_542
timestamp 1675432918
transform 1 0 12650 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_543
timestamp 1675432918
transform 1 0 12650 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_544
timestamp 1675432918
transform 1 0 12650 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_545
timestamp 1675432918
transform 1 0 12650 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_546
timestamp 1675432918
transform 1 0 12650 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_547
timestamp 1675432918
transform 1 0 12650 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_548
timestamp 1675432918
transform 1 0 12650 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_549
timestamp 1675432918
transform 1 0 12650 0 1 22550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_550
timestamp 1675432918
transform 1 0 12650 0 1 23650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_551
timestamp 1675432918
transform 1 0 12650 0 1 24750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_552
timestamp 1675432918
transform 1 0 13200 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_553
timestamp 1675432918
transform 1 0 13200 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_554
timestamp 1675432918
transform 1 0 13200 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_555
timestamp 1675432918
transform 1 0 13200 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_556
timestamp 1675432918
transform 1 0 13200 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_557
timestamp 1675432918
transform 1 0 13200 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_558
timestamp 1675432918
transform 1 0 13200 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_559
timestamp 1675432918
transform 1 0 13200 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_560
timestamp 1675432918
transform 1 0 13200 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_561
timestamp 1675432918
transform 1 0 13200 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_562
timestamp 1675432918
transform 1 0 13200 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_563
timestamp 1675432918
transform 1 0 13200 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_564
timestamp 1675432918
transform 1 0 13200 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_565
timestamp 1675432918
transform 1 0 13200 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_566
timestamp 1675432918
transform 1 0 13200 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_567
timestamp 1675432918
transform 1 0 13200 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_568
timestamp 1675432918
transform 1 0 13200 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_569
timestamp 1675432918
transform 1 0 13200 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_570
timestamp 1675432918
transform 1 0 13200 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_571
timestamp 1675432918
transform 1 0 13200 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_572
timestamp 1675432918
transform 1 0 13200 0 1 22000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_573
timestamp 1675432918
transform 1 0 13200 0 1 23100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_574
timestamp 1675432918
transform 1 0 13200 0 1 24200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_575
timestamp 1675432918
transform 1 0 13750 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_576
timestamp 1675432918
transform 1 0 13750 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_577
timestamp 1675432918
transform 1 0 13750 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_578
timestamp 1675432918
transform 1 0 13750 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_579
timestamp 1675432918
transform 1 0 13750 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_580
timestamp 1675432918
transform 1 0 13750 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_581
timestamp 1675432918
transform 1 0 13750 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_582
timestamp 1675432918
transform 1 0 13750 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_583
timestamp 1675432918
transform 1 0 13750 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_584
timestamp 1675432918
transform 1 0 13750 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_585
timestamp 1675432918
transform 1 0 13750 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_586
timestamp 1675432918
transform 1 0 13750 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_587
timestamp 1675432918
transform 1 0 13750 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_588
timestamp 1675432918
transform 1 0 13750 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_589
timestamp 1675432918
transform 1 0 13750 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_590
timestamp 1675432918
transform 1 0 13750 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_591
timestamp 1675432918
transform 1 0 13750 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_592
timestamp 1675432918
transform 1 0 13750 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_593
timestamp 1675432918
transform 1 0 13750 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_594
timestamp 1675432918
transform 1 0 13750 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_595
timestamp 1675432918
transform 1 0 13750 0 1 22550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_596
timestamp 1675432918
transform 1 0 13750 0 1 23650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_597
timestamp 1675432918
transform 1 0 13750 0 1 24750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_598
timestamp 1675432918
transform 1 0 14300 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_599
timestamp 1675432918
transform 1 0 14300 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_600
timestamp 1675432918
transform 1 0 14300 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_601
timestamp 1675432918
transform 1 0 14300 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_602
timestamp 1675432918
transform 1 0 14300 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_603
timestamp 1675432918
transform 1 0 14300 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_604
timestamp 1675432918
transform 1 0 14300 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_605
timestamp 1675432918
transform 1 0 14300 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_606
timestamp 1675432918
transform 1 0 14300 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_607
timestamp 1675432918
transform 1 0 14300 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_608
timestamp 1675432918
transform 1 0 14300 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_609
timestamp 1675432918
transform 1 0 14300 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_610
timestamp 1675432918
transform 1 0 14300 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_611
timestamp 1675432918
transform 1 0 14300 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_612
timestamp 1675432918
transform 1 0 14300 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_613
timestamp 1675432918
transform 1 0 14300 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_614
timestamp 1675432918
transform 1 0 14300 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_615
timestamp 1675432918
transform 1 0 14300 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_616
timestamp 1675432918
transform 1 0 14300 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_617
timestamp 1675432918
transform 1 0 14300 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_618
timestamp 1675432918
transform 1 0 14300 0 1 22000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_619
timestamp 1675432918
transform 1 0 14300 0 1 23100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_620
timestamp 1675432918
transform 1 0 14300 0 1 24200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_621
timestamp 1675432918
transform 1 0 14850 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_622
timestamp 1675432918
transform 1 0 14850 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_623
timestamp 1675432918
transform 1 0 14850 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_624
timestamp 1675432918
transform 1 0 14850 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_625
timestamp 1675432918
transform 1 0 14850 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_626
timestamp 1675432918
transform 1 0 14850 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_627
timestamp 1675432918
transform 1 0 14850 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_628
timestamp 1675432918
transform 1 0 14850 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_629
timestamp 1675432918
transform 1 0 14850 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_630
timestamp 1675432918
transform 1 0 14850 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_631
timestamp 1675432918
transform 1 0 14850 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_632
timestamp 1675432918
transform 1 0 14850 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_633
timestamp 1675432918
transform 1 0 14850 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_634
timestamp 1675432918
transform 1 0 14850 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_635
timestamp 1675432918
transform 1 0 14850 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_636
timestamp 1675432918
transform 1 0 14850 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_637
timestamp 1675432918
transform 1 0 14850 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_638
timestamp 1675432918
transform 1 0 14850 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_639
timestamp 1675432918
transform 1 0 14850 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_640
timestamp 1675432918
transform 1 0 14850 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_641
timestamp 1675432918
transform 1 0 14850 0 1 22550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_642
timestamp 1675432918
transform 1 0 14850 0 1 23650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_643
timestamp 1675432918
transform 1 0 14850 0 1 24750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_644
timestamp 1675432918
transform 1 0 15400 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_645
timestamp 1675432918
transform 1 0 15400 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_646
timestamp 1675432918
transform 1 0 15400 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_647
timestamp 1675432918
transform 1 0 15400 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_648
timestamp 1675432918
transform 1 0 15400 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_649
timestamp 1675432918
transform 1 0 15400 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_650
timestamp 1675432918
transform 1 0 15400 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_651
timestamp 1675432918
transform 1 0 15400 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_652
timestamp 1675432918
transform 1 0 15400 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_653
timestamp 1675432918
transform 1 0 15400 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_654
timestamp 1675432918
transform 1 0 15400 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_655
timestamp 1675432918
transform 1 0 15400 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_656
timestamp 1675432918
transform 1 0 15400 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_657
timestamp 1675432918
transform 1 0 15400 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_658
timestamp 1675432918
transform 1 0 15400 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_659
timestamp 1675432918
transform 1 0 15400 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_660
timestamp 1675432918
transform 1 0 15400 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_661
timestamp 1675432918
transform 1 0 15400 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_662
timestamp 1675432918
transform 1 0 15400 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_663
timestamp 1675432918
transform 1 0 15400 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_664
timestamp 1675432918
transform 1 0 15400 0 1 22000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_665
timestamp 1675432918
transform 1 0 15400 0 1 23100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_666
timestamp 1675432918
transform 1 0 15400 0 1 24200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_667
timestamp 1675432918
transform 1 0 15950 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_668
timestamp 1675432918
transform 1 0 15950 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_669
timestamp 1675432918
transform 1 0 15950 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_670
timestamp 1675432918
transform 1 0 15950 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_671
timestamp 1675432918
transform 1 0 15950 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_672
timestamp 1675432918
transform 1 0 15950 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_673
timestamp 1675432918
transform 1 0 15950 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_674
timestamp 1675432918
transform 1 0 15950 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_675
timestamp 1675432918
transform 1 0 15950 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_676
timestamp 1675432918
transform 1 0 15950 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_677
timestamp 1675432918
transform 1 0 15950 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_678
timestamp 1675432918
transform 1 0 15950 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_679
timestamp 1675432918
transform 1 0 15950 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_680
timestamp 1675432918
transform 1 0 15950 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_681
timestamp 1675432918
transform 1 0 15950 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_682
timestamp 1675432918
transform 1 0 15950 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_683
timestamp 1675432918
transform 1 0 15950 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_684
timestamp 1675432918
transform 1 0 15950 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_685
timestamp 1675432918
transform 1 0 15950 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_686
timestamp 1675432918
transform 1 0 15950 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_687
timestamp 1675432918
transform 1 0 15950 0 1 22550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_688
timestamp 1675432918
transform 1 0 15950 0 1 23650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_689
timestamp 1675432918
transform 1 0 15950 0 1 24750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_690
timestamp 1675432918
transform 1 0 16500 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_691
timestamp 1675432918
transform 1 0 16500 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_692
timestamp 1675432918
transform 1 0 16500 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_693
timestamp 1675432918
transform 1 0 16500 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_694
timestamp 1675432918
transform 1 0 16500 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_695
timestamp 1675432918
transform 1 0 16500 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_696
timestamp 1675432918
transform 1 0 16500 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_697
timestamp 1675432918
transform 1 0 16500 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_698
timestamp 1675432918
transform 1 0 16500 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_699
timestamp 1675432918
transform 1 0 16500 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_700
timestamp 1675432918
transform 1 0 16500 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_701
timestamp 1675432918
transform 1 0 16500 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_702
timestamp 1675432918
transform 1 0 16500 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_703
timestamp 1675432918
transform 1 0 16500 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_704
timestamp 1675432918
transform 1 0 16500 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_705
timestamp 1675432918
transform 1 0 16500 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_706
timestamp 1675432918
transform 1 0 16500 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_707
timestamp 1675432918
transform 1 0 16500 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_708
timestamp 1675432918
transform 1 0 16500 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_709
timestamp 1675432918
transform 1 0 16500 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_710
timestamp 1675432918
transform 1 0 16500 0 1 22000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_711
timestamp 1675432918
transform 1 0 16500 0 1 23100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_712
timestamp 1675432918
transform 1 0 16500 0 1 24200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_713
timestamp 1675432918
transform 1 0 17050 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_714
timestamp 1675432918
transform 1 0 17050 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_715
timestamp 1675432918
transform 1 0 17050 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_716
timestamp 1675432918
transform 1 0 17050 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_717
timestamp 1675432918
transform 1 0 17050 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_718
timestamp 1675432918
transform 1 0 17050 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_719
timestamp 1675432918
transform 1 0 17050 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_720
timestamp 1675432918
transform 1 0 17050 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_721
timestamp 1675432918
transform 1 0 17050 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_722
timestamp 1675432918
transform 1 0 17050 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_723
timestamp 1675432918
transform 1 0 17050 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_724
timestamp 1675432918
transform 1 0 17050 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_725
timestamp 1675432918
transform 1 0 17050 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_726
timestamp 1675432918
transform 1 0 17050 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_727
timestamp 1675432918
transform 1 0 17050 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_728
timestamp 1675432918
transform 1 0 17050 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_729
timestamp 1675432918
transform 1 0 17050 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_730
timestamp 1675432918
transform 1 0 17050 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_731
timestamp 1675432918
transform 1 0 17050 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_732
timestamp 1675432918
transform 1 0 17050 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_733
timestamp 1675432918
transform 1 0 17050 0 1 22550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_734
timestamp 1675432918
transform 1 0 17050 0 1 23650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_735
timestamp 1675432918
transform 1 0 17050 0 1 24750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_736
timestamp 1675432918
transform 1 0 17600 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_737
timestamp 1675432918
transform 1 0 17600 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_738
timestamp 1675432918
transform 1 0 17600 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_739
timestamp 1675432918
transform 1 0 17600 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_740
timestamp 1675432918
transform 1 0 17600 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_741
timestamp 1675432918
transform 1 0 17600 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_742
timestamp 1675432918
transform 1 0 17600 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_743
timestamp 1675432918
transform 1 0 17600 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_744
timestamp 1675432918
transform 1 0 17600 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_745
timestamp 1675432918
transform 1 0 17600 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_746
timestamp 1675432918
transform 1 0 17600 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_747
timestamp 1675432918
transform 1 0 17600 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_748
timestamp 1675432918
transform 1 0 17600 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_749
timestamp 1675432918
transform 1 0 17600 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_750
timestamp 1675432918
transform 1 0 17600 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_751
timestamp 1675432918
transform 1 0 17600 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_752
timestamp 1675432918
transform 1 0 17600 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_753
timestamp 1675432918
transform 1 0 17600 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_754
timestamp 1675432918
transform 1 0 17600 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_755
timestamp 1675432918
transform 1 0 17600 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_756
timestamp 1675432918
transform 1 0 17600 0 1 22000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_757
timestamp 1675432918
transform 1 0 17600 0 1 23100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_758
timestamp 1675432918
transform 1 0 17600 0 1 24200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_759
timestamp 1675432918
transform 1 0 18150 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_760
timestamp 1675432918
transform 1 0 18150 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_761
timestamp 1675432918
transform 1 0 18150 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_762
timestamp 1675432918
transform 1 0 18150 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_763
timestamp 1675432918
transform 1 0 18150 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_764
timestamp 1675432918
transform 1 0 18150 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_765
timestamp 1675432918
transform 1 0 18150 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_766
timestamp 1675432918
transform 1 0 18150 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_767
timestamp 1675432918
transform 1 0 18150 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_768
timestamp 1675432918
transform 1 0 18150 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_769
timestamp 1675432918
transform 1 0 18150 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_770
timestamp 1675432918
transform 1 0 18150 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_771
timestamp 1675432918
transform 1 0 18150 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_772
timestamp 1675432918
transform 1 0 18150 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_773
timestamp 1675432918
transform 1 0 18150 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_774
timestamp 1675432918
transform 1 0 18150 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_775
timestamp 1675432918
transform 1 0 18150 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_776
timestamp 1675432918
transform 1 0 18150 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_777
timestamp 1675432918
transform 1 0 18150 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_778
timestamp 1675432918
transform 1 0 18150 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_779
timestamp 1675432918
transform 1 0 18150 0 1 22550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_780
timestamp 1675432918
transform 1 0 18150 0 1 23650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_781
timestamp 1675432918
transform 1 0 18150 0 1 24750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_782
timestamp 1675432918
transform 1 0 18700 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_783
timestamp 1675432918
transform 1 0 18700 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_784
timestamp 1675432918
transform 1 0 18700 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_785
timestamp 1675432918
transform 1 0 18700 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_786
timestamp 1675432918
transform 1 0 18700 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_787
timestamp 1675432918
transform 1 0 18700 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_788
timestamp 1675432918
transform 1 0 18700 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_789
timestamp 1675432918
transform 1 0 18700 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_790
timestamp 1675432918
transform 1 0 18700 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_791
timestamp 1675432918
transform 1 0 18700 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_792
timestamp 1675432918
transform 1 0 18700 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_793
timestamp 1675432918
transform 1 0 18700 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_794
timestamp 1675432918
transform 1 0 18700 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_795
timestamp 1675432918
transform 1 0 18700 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_796
timestamp 1675432918
transform 1 0 18700 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_797
timestamp 1675432918
transform 1 0 18700 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_798
timestamp 1675432918
transform 1 0 18700 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_799
timestamp 1675432918
transform 1 0 18700 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_800
timestamp 1675432918
transform 1 0 18700 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_801
timestamp 1675432918
transform 1 0 18700 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_802
timestamp 1675432918
transform 1 0 18700 0 1 22000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_803
timestamp 1675432918
transform 1 0 18700 0 1 23100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_804
timestamp 1675432918
transform 1 0 18700 0 1 24200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_805
timestamp 1675432918
transform 1 0 19250 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_806
timestamp 1675432918
transform 1 0 19250 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_807
timestamp 1675432918
transform 1 0 19250 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_808
timestamp 1675432918
transform 1 0 19250 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_809
timestamp 1675432918
transform 1 0 19250 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_810
timestamp 1675432918
transform 1 0 19250 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_811
timestamp 1675432918
transform 1 0 19250 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_812
timestamp 1675432918
transform 1 0 19250 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_813
timestamp 1675432918
transform 1 0 19250 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_814
timestamp 1675432918
transform 1 0 19250 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_815
timestamp 1675432918
transform 1 0 19250 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_816
timestamp 1675432918
transform 1 0 19250 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_817
timestamp 1675432918
transform 1 0 19250 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_818
timestamp 1675432918
transform 1 0 19250 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_819
timestamp 1675432918
transform 1 0 19250 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_820
timestamp 1675432918
transform 1 0 19250 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_821
timestamp 1675432918
transform 1 0 19250 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_822
timestamp 1675432918
transform 1 0 19250 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_823
timestamp 1675432918
transform 1 0 19250 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_824
timestamp 1675432918
transform 1 0 19250 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_825
timestamp 1675432918
transform 1 0 19250 0 1 22550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_826
timestamp 1675432918
transform 1 0 19250 0 1 23650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_827
timestamp 1675432918
transform 1 0 19250 0 1 24750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_828
timestamp 1675432918
transform 1 0 19800 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_829
timestamp 1675432918
transform 1 0 19800 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_830
timestamp 1675432918
transform 1 0 19800 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_831
timestamp 1675432918
transform 1 0 19800 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_832
timestamp 1675432918
transform 1 0 19800 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_833
timestamp 1675432918
transform 1 0 19800 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_834
timestamp 1675432918
transform 1 0 19800 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_835
timestamp 1675432918
transform 1 0 19800 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_836
timestamp 1675432918
transform 1 0 19800 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_837
timestamp 1675432918
transform 1 0 19800 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_838
timestamp 1675432918
transform 1 0 19800 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_839
timestamp 1675432918
transform 1 0 19800 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_840
timestamp 1675432918
transform 1 0 19800 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_841
timestamp 1675432918
transform 1 0 19800 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_842
timestamp 1675432918
transform 1 0 19800 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_843
timestamp 1675432918
transform 1 0 19800 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_844
timestamp 1675432918
transform 1 0 19800 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_845
timestamp 1675432918
transform 1 0 19800 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_846
timestamp 1675432918
transform 1 0 19800 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_847
timestamp 1675432918
transform 1 0 19800 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_848
timestamp 1675432918
transform 1 0 19800 0 1 22000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_849
timestamp 1675432918
transform 1 0 19800 0 1 23100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_850
timestamp 1675432918
transform 1 0 19800 0 1 24200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_851
timestamp 1675432918
transform 1 0 20350 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_852
timestamp 1675432918
transform 1 0 20350 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_853
timestamp 1675432918
transform 1 0 20350 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_854
timestamp 1675432918
transform 1 0 20350 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_855
timestamp 1675432918
transform 1 0 20350 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_856
timestamp 1675432918
transform 1 0 20350 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_857
timestamp 1675432918
transform 1 0 20350 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_858
timestamp 1675432918
transform 1 0 20350 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_859
timestamp 1675432918
transform 1 0 20350 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_860
timestamp 1675432918
transform 1 0 20350 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_861
timestamp 1675432918
transform 1 0 20350 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_862
timestamp 1675432918
transform 1 0 20350 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_863
timestamp 1675432918
transform 1 0 20350 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_864
timestamp 1675432918
transform 1 0 20350 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_865
timestamp 1675432918
transform 1 0 20350 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_866
timestamp 1675432918
transform 1 0 20350 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_867
timestamp 1675432918
transform 1 0 20350 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_868
timestamp 1675432918
transform 1 0 20350 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_869
timestamp 1675432918
transform 1 0 20350 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_870
timestamp 1675432918
transform 1 0 20350 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_871
timestamp 1675432918
transform 1 0 20350 0 1 22550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_872
timestamp 1675432918
transform 1 0 20350 0 1 23650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_873
timestamp 1675432918
transform 1 0 20350 0 1 24750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_874
timestamp 1675432918
transform 1 0 20900 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_875
timestamp 1675432918
transform 1 0 20900 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_876
timestamp 1675432918
transform 1 0 20900 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_877
timestamp 1675432918
transform 1 0 20900 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_878
timestamp 1675432918
transform 1 0 20900 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_879
timestamp 1675432918
transform 1 0 20900 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_880
timestamp 1675432918
transform 1 0 20900 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_881
timestamp 1675432918
transform 1 0 20900 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_882
timestamp 1675432918
transform 1 0 20900 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_883
timestamp 1675432918
transform 1 0 20900 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_884
timestamp 1675432918
transform 1 0 20900 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_885
timestamp 1675432918
transform 1 0 20900 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_886
timestamp 1675432918
transform 1 0 20900 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_887
timestamp 1675432918
transform 1 0 20900 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_888
timestamp 1675432918
transform 1 0 20900 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_889
timestamp 1675432918
transform 1 0 20900 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_890
timestamp 1675432918
transform 1 0 20900 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_891
timestamp 1675432918
transform 1 0 20900 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_892
timestamp 1675432918
transform 1 0 20900 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_893
timestamp 1675432918
transform 1 0 20900 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_894
timestamp 1675432918
transform 1 0 20900 0 1 22000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_895
timestamp 1675432918
transform 1 0 20900 0 1 23100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_896
timestamp 1675432918
transform 1 0 20900 0 1 24200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_897
timestamp 1675432918
transform 1 0 21450 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_898
timestamp 1675432918
transform 1 0 21450 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_899
timestamp 1675432918
transform 1 0 21450 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_900
timestamp 1675432918
transform 1 0 21450 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_901
timestamp 1675432918
transform 1 0 21450 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_902
timestamp 1675432918
transform 1 0 21450 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_903
timestamp 1675432918
transform 1 0 21450 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_904
timestamp 1675432918
transform 1 0 21450 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_905
timestamp 1675432918
transform 1 0 21450 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_906
timestamp 1675432918
transform 1 0 21450 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_907
timestamp 1675432918
transform 1 0 21450 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_908
timestamp 1675432918
transform 1 0 21450 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_909
timestamp 1675432918
transform 1 0 21450 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_910
timestamp 1675432918
transform 1 0 21450 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_911
timestamp 1675432918
transform 1 0 21450 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_912
timestamp 1675432918
transform 1 0 21450 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_913
timestamp 1675432918
transform 1 0 21450 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_914
timestamp 1675432918
transform 1 0 21450 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_915
timestamp 1675432918
transform 1 0 21450 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_916
timestamp 1675432918
transform 1 0 21450 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_917
timestamp 1675432918
transform 1 0 21450 0 1 22550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_918
timestamp 1675432918
transform 1 0 21450 0 1 23650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_919
timestamp 1675432918
transform 1 0 21450 0 1 24750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_920
timestamp 1675432918
transform 1 0 22000 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_921
timestamp 1675432918
transform 1 0 22000 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_922
timestamp 1675432918
transform 1 0 22000 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_923
timestamp 1675432918
transform 1 0 22000 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_924
timestamp 1675432918
transform 1 0 22000 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_925
timestamp 1675432918
transform 1 0 22000 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_926
timestamp 1675432918
transform 1 0 22000 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_927
timestamp 1675432918
transform 1 0 22000 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_928
timestamp 1675432918
transform 1 0 22000 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_929
timestamp 1675432918
transform 1 0 22000 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_930
timestamp 1675432918
transform 1 0 22000 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_931
timestamp 1675432918
transform 1 0 22000 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_932
timestamp 1675432918
transform 1 0 22000 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_933
timestamp 1675432918
transform 1 0 22000 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_934
timestamp 1675432918
transform 1 0 22000 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_935
timestamp 1675432918
transform 1 0 22000 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_936
timestamp 1675432918
transform 1 0 22000 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_937
timestamp 1675432918
transform 1 0 22000 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_938
timestamp 1675432918
transform 1 0 22000 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_939
timestamp 1675432918
transform 1 0 22000 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_940
timestamp 1675432918
transform 1 0 22000 0 1 22000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_941
timestamp 1675432918
transform 1 0 22000 0 1 23100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_942
timestamp 1675432918
transform 1 0 22000 0 1 24200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_943
timestamp 1675432918
transform 1 0 22550 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_944
timestamp 1675432918
transform 1 0 22550 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_945
timestamp 1675432918
transform 1 0 22550 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_946
timestamp 1675432918
transform 1 0 22550 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_947
timestamp 1675432918
transform 1 0 22550 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_948
timestamp 1675432918
transform 1 0 22550 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_949
timestamp 1675432918
transform 1 0 22550 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_950
timestamp 1675432918
transform 1 0 22550 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_951
timestamp 1675432918
transform 1 0 22550 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_952
timestamp 1675432918
transform 1 0 22550 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_953
timestamp 1675432918
transform 1 0 22550 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_954
timestamp 1675432918
transform 1 0 22550 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_955
timestamp 1675432918
transform 1 0 22550 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_956
timestamp 1675432918
transform 1 0 22550 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_957
timestamp 1675432918
transform 1 0 22550 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_958
timestamp 1675432918
transform 1 0 22550 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_959
timestamp 1675432918
transform 1 0 22550 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_960
timestamp 1675432918
transform 1 0 22550 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_961
timestamp 1675432918
transform 1 0 22550 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_962
timestamp 1675432918
transform 1 0 22550 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_963
timestamp 1675432918
transform 1 0 22550 0 1 22550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_964
timestamp 1675432918
transform 1 0 22550 0 1 23650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_965
timestamp 1675432918
transform 1 0 22550 0 1 24750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_966
timestamp 1675432918
transform 1 0 23100 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_967
timestamp 1675432918
transform 1 0 23100 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_968
timestamp 1675432918
transform 1 0 23100 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_969
timestamp 1675432918
transform 1 0 23100 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_970
timestamp 1675432918
transform 1 0 23100 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_971
timestamp 1675432918
transform 1 0 23100 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_972
timestamp 1675432918
transform 1 0 23100 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_973
timestamp 1675432918
transform 1 0 23100 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_974
timestamp 1675432918
transform 1 0 23100 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_975
timestamp 1675432918
transform 1 0 23100 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_976
timestamp 1675432918
transform 1 0 23100 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_977
timestamp 1675432918
transform 1 0 23100 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_978
timestamp 1675432918
transform 1 0 23100 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_979
timestamp 1675432918
transform 1 0 23100 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_980
timestamp 1675432918
transform 1 0 23100 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_981
timestamp 1675432918
transform 1 0 23100 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_982
timestamp 1675432918
transform 1 0 23100 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_983
timestamp 1675432918
transform 1 0 23100 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_984
timestamp 1675432918
transform 1 0 23100 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_985
timestamp 1675432918
transform 1 0 23100 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_986
timestamp 1675432918
transform 1 0 23100 0 1 22000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_987
timestamp 1675432918
transform 1 0 23100 0 1 23100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_988
timestamp 1675432918
transform 1 0 23100 0 1 24200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_989
timestamp 1675432918
transform 1 0 23650 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_990
timestamp 1675432918
transform 1 0 23650 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_991
timestamp 1675432918
transform 1 0 23650 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_992
timestamp 1675432918
transform 1 0 23650 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_993
timestamp 1675432918
transform 1 0 23650 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_994
timestamp 1675432918
transform 1 0 23650 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_995
timestamp 1675432918
transform 1 0 23650 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_996
timestamp 1675432918
transform 1 0 23650 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_997
timestamp 1675432918
transform 1 0 23650 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_998
timestamp 1675432918
transform 1 0 23650 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_999
timestamp 1675432918
transform 1 0 23650 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1000
timestamp 1675432918
transform 1 0 23650 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1001
timestamp 1675432918
transform 1 0 23650 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1002
timestamp 1675432918
transform 1 0 23650 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1003
timestamp 1675432918
transform 1 0 23650 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1004
timestamp 1675432918
transform 1 0 23650 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1005
timestamp 1675432918
transform 1 0 23650 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1006
timestamp 1675432918
transform 1 0 23650 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1007
timestamp 1675432918
transform 1 0 23650 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1008
timestamp 1675432918
transform 1 0 23650 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1009
timestamp 1675432918
transform 1 0 23650 0 1 22550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1010
timestamp 1675432918
transform 1 0 23650 0 1 23650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1011
timestamp 1675432918
transform 1 0 23650 0 1 24750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1012
timestamp 1675432918
transform 1 0 24200 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1013
timestamp 1675432918
transform 1 0 24200 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1014
timestamp 1675432918
transform 1 0 24200 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1015
timestamp 1675432918
transform 1 0 24200 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1016
timestamp 1675432918
transform 1 0 24200 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1017
timestamp 1675432918
transform 1 0 24200 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1018
timestamp 1675432918
transform 1 0 24200 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1019
timestamp 1675432918
transform 1 0 24200 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1020
timestamp 1675432918
transform 1 0 24200 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1021
timestamp 1675432918
transform 1 0 24200 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1022
timestamp 1675432918
transform 1 0 24200 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1023
timestamp 1675432918
transform 1 0 24200 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1024
timestamp 1675432918
transform 1 0 24200 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1025
timestamp 1675432918
transform 1 0 24200 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1026
timestamp 1675432918
transform 1 0 24200 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1027
timestamp 1675432918
transform 1 0 24200 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1028
timestamp 1675432918
transform 1 0 24200 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1029
timestamp 1675432918
transform 1 0 24200 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1030
timestamp 1675432918
transform 1 0 24200 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1031
timestamp 1675432918
transform 1 0 24200 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1032
timestamp 1675432918
transform 1 0 24200 0 1 22000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1033
timestamp 1675432918
transform 1 0 24200 0 1 23100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1034
timestamp 1675432918
transform 1 0 24200 0 1 24200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1035
timestamp 1675432918
transform 1 0 24750 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1036
timestamp 1675432918
transform 1 0 24750 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1037
timestamp 1675432918
transform 1 0 24750 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1038
timestamp 1675432918
transform 1 0 24750 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1039
timestamp 1675432918
transform 1 0 24750 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1040
timestamp 1675432918
transform 1 0 24750 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1041
timestamp 1675432918
transform 1 0 24750 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1042
timestamp 1675432918
transform 1 0 24750 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1043
timestamp 1675432918
transform 1 0 24750 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1044
timestamp 1675432918
transform 1 0 24750 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1045
timestamp 1675432918
transform 1 0 24750 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1046
timestamp 1675432918
transform 1 0 24750 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1047
timestamp 1675432918
transform 1 0 24750 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1048
timestamp 1675432918
transform 1 0 24750 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1049
timestamp 1675432918
transform 1 0 24750 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1050
timestamp 1675432918
transform 1 0 24750 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1051
timestamp 1675432918
transform 1 0 24750 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1052
timestamp 1675432918
transform 1 0 24750 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1053
timestamp 1675432918
transform 1 0 24750 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1054
timestamp 1675432918
transform 1 0 24750 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1055
timestamp 1675432918
transform 1 0 24750 0 1 22550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1056
timestamp 1675432918
transform 1 0 24750 0 1 23650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1057
timestamp 1675432918
transform 1 0 24750 0 1 24750
box -113 -113 663 663
<< end >>
