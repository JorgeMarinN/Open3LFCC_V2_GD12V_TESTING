magic
tech sky130A
timestamp 1699898483
<< metal2 >>
rect 3000 56640 6800 58000
rect 3000 56400 5740 56640
rect 5930 56400 6800 56640
rect 3000 5749 4962 6000
rect 3000 5200 5300 5749
<< metal3 >>
rect 6000 58000 30000 61000
rect 1000 35000 4000 56000
rect 27000 37000 30000 58000
rect 1000 27000 25000 35000
rect 1000 7000 4000 27000
rect 27000 4000 30000 25000
rect 6000 1000 30000 4000
<< metal4 >>
rect 6000 58000 30000 61000
rect 1000 35000 4000 56000
rect 27000 37000 30000 58000
rect 1000 27000 25000 35000
rect 1000 7000 4000 27000
rect 27000 4000 30000 25000
rect 6000 1000 30000 4000
<< metal5 >>
rect 6000 58000 30000 61000
rect 1000 35000 4000 56000
rect 27000 37000 30000 58000
rect 1000 27000 25000 35000
rect 1000 7000 4000 27000
rect 27000 4000 30000 25000
rect 6000 1000 30000 4000
use nmos_waffle_36x36  nmos_waffle_36x36_0
timestamp 1693601174
transform 1 0 5925 0 1 5975
box -5925 -5975 24675 24625
use nmos_waffle_36x36  nmos_waffle_36x36_1
timestamp 1693601174
transform 0 1 5975 -1 0 55675
box -5925 -5975 24675 24625
<< labels >>
rlabel metal5 6000 58900 7000 59900 7 VP
rlabel metal5 2000 30500 6000 31500 7 out
rlabel metal5 6000 2000 7000 3000 7 VN
rlabel metal2 3000 57000 4000 58000 7 s2
rlabel metal2 3000 5500 4000 6000 7 s1
rlabel space 2881 2944 2881 2944 7 DNW1
rlabel space 2881 59700 2881 59700 7 DNW2
<< end >>
