magic
tech sky130A
magscale 1 2
timestamp 1700232449
<< nwell >>
rect 682 261 740 582
<< pwell >>
rect 760 885 1680 1067
rect 3 38 3018 204
<< locali >>
rect 777 1020 835 1100
rect 680 828 980 872
rect 1020 828 1200 872
rect 17 460 75 540
rect 220 215 480 263
rect 680 257 720 828
rect 777 460 835 620
rect 540 256 720 257
rect 540 222 680 256
rect 714 222 720 256
rect 1960 254 2160 262
rect 540 215 720 222
rect 1960 220 2040 254
rect 2074 220 2160 254
rect 2200 220 2400 262
rect 17 0 75 100
rect 777 0 835 100
rect 260 -114 340 -100
rect 260 -166 274 -114
rect 326 -166 340 -114
rect 260 -180 340 -166
rect 3040 -114 3120 -100
rect 3040 -166 3054 -114
rect 3106 -166 3120 -114
rect 3040 -180 3120 -166
rect 263 -560 305 -180
rect 3055 -560 3097 -180
<< viali >>
rect 1344 838 1378 872
rect 1526 840 1560 874
rect 126 215 160 249
rect 680 222 714 256
rect 1000 222 1100 256
rect 1620 220 1654 254
rect 1840 220 1874 254
rect 2040 220 2074 254
rect 2520 220 2554 254
rect 2706 220 2740 260
rect 274 -166 326 -114
rect 3054 -166 3106 -114
<< metal1 >>
rect 3260 1136 3360 1140
rect 0 1040 3360 1136
rect 1324 888 1404 898
rect 1324 828 1334 888
rect 1394 828 1404 888
rect 1324 818 1404 828
rect 1506 874 1580 894
rect 1506 840 1526 874
rect 1560 840 1580 874
rect 1506 820 1580 840
rect 0 572 3020 592
rect 0 512 140 572
rect 200 512 3020 572
rect 0 496 3020 512
rect 1090 358 2560 412
rect 1090 280 1136 358
rect 2520 280 2560 358
rect 0 249 200 280
rect 0 215 126 249
rect 160 215 200 249
rect 0 200 200 215
rect 660 260 734 280
rect 980 260 1136 280
rect 660 256 1136 260
rect 660 222 680 256
rect 714 222 1000 256
rect 1100 222 1136 256
rect 660 220 1136 222
rect 660 200 734 220
rect 980 200 1136 220
rect 1600 270 1680 280
rect 1600 210 1610 270
rect 1670 210 1680 270
rect 1600 200 1680 210
rect 1820 270 1900 280
rect 1820 210 1830 270
rect 1890 210 1900 270
rect 1820 200 1900 210
rect 2020 270 2100 280
rect 2020 210 2030 270
rect 2090 210 2100 270
rect 2020 200 2100 210
rect 2500 254 2580 280
rect 2500 220 2520 254
rect 2554 220 2580 254
rect 2500 200 2580 220
rect 2680 260 2760 280
rect 2680 220 2706 260
rect 2740 220 2760 260
rect 2680 200 2760 220
rect 1090 198 1136 200
rect 2520 192 2560 200
rect 0 -48 3020 48
rect 3260 -60 3360 1040
rect 260 -114 340 -100
rect 260 -166 274 -114
rect 326 -166 340 -114
rect 260 -180 340 -166
rect 3040 -114 3120 -100
rect 3040 -166 3054 -114
rect 3106 -166 3120 -114
rect 3040 -180 3120 -166
<< via1 >>
rect 1334 872 1394 888
rect 1334 838 1344 872
rect 1344 838 1378 872
rect 1378 838 1394 872
rect 1334 828 1394 838
rect 140 512 200 572
rect 1610 254 1670 270
rect 1610 220 1620 254
rect 1620 220 1654 254
rect 1654 220 1670 254
rect 1610 210 1670 220
rect 1830 254 1890 270
rect 1830 220 1840 254
rect 1840 220 1874 254
rect 1874 220 1890 254
rect 1830 210 1890 220
rect 2030 254 2090 270
rect 2030 220 2040 254
rect 2040 220 2074 254
rect 2074 220 2090 254
rect 2030 210 2090 220
rect 274 -166 326 -114
rect 3054 -166 3106 -114
rect 564 -380 620 -320
rect 1652 -380 1708 -320
rect 2740 -380 2796 -320
<< metal2 >>
rect 1304 888 1418 912
rect 1304 828 1334 888
rect 1394 828 1418 888
rect 1304 800 1418 828
rect 1340 700 1380 800
rect 1340 660 2080 700
rect 120 572 220 592
rect 120 512 140 572
rect 200 512 220 572
rect 120 -300 220 512
rect 2040 300 2080 660
rect 1580 270 1700 300
rect 1580 210 1610 270
rect 1670 210 1700 270
rect 1580 180 1700 210
rect 1800 270 1920 300
rect 1800 210 1830 270
rect 1890 210 1920 270
rect 1800 180 1920 210
rect 2000 270 2120 300
rect 2000 210 2030 270
rect 2090 210 2120 270
rect 2000 180 2120 210
rect 1600 -100 1660 180
rect 260 -114 1660 -100
rect 260 -166 274 -114
rect 326 -160 1660 -114
rect 1820 -100 1880 180
rect 1820 -114 3120 -100
rect 1820 -160 3054 -114
rect 326 -166 340 -160
rect 260 -180 340 -166
rect 3040 -166 3054 -160
rect 3106 -166 3120 -114
rect 3040 -180 3120 -166
rect 120 -320 2816 -300
rect 120 -380 564 -320
rect 620 -380 1652 -320
rect 1708 -380 2740 -320
rect 2796 -380 2816 -320
rect 120 -400 2816 -380
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 2308 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_1
timestamp 1683767628
transform 1 0 1128 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 368 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1683767628
transform 1 0 1756 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1683767628
transform 1 0 2032 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1683767628
transform 1 0 852 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 92 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  sky130_fd_sc_hd__inv_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 852 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 0 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_1
timestamp 1683767628
transform 1 0 760 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_2
timestamp 1683767628
transform 1 0 760 0 -1 1088
box -38 -48 130 592
use sp_delay_top  sp_delay_top_0
timestamp 1700231096
transform 0 1 0 -1 0 42
box 0 0 6422 3360
<< labels >>
rlabel metal1 3260 1040 3360 1140 1 VSS
port 1 n
rlabel metal2 120 492 220 592 1 VCC
port 2 n
rlabel metal1 0 200 80 280 7 Vin
port 3 w
rlabel metal1 1506 820 1580 894 3 VFE
port 4 e
rlabel metal1 2680 200 2760 280 3 VRE
port 5 e
<< end >>
