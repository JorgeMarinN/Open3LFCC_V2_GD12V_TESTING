magic
tech sky130A
magscale 1 2
timestamp 1699972156
<< pwell >>
rect -53 -53 2763 2763
<< psubdiff >>
rect -17 2693 79 2727
rect 2631 2693 2727 2727
rect -17 17 17 2693
rect 2693 2631 2727 2693
rect 2693 17 2727 79
rect -17 -17 79 17
rect 2631 -17 2727 17
<< psubdiffcont >>
rect 79 2693 2631 2727
rect 2693 79 2727 2631
rect 79 -17 2631 17
<< ndiode >>
rect 85 2613 2625 2625
rect 85 97 97 2613
rect 2613 97 2625 2613
rect 85 85 2625 97
<< ndiodec >>
rect 97 97 2613 2613
<< locali >>
rect -17 2693 79 2727
rect 2631 2693 2727 2727
rect -17 17 17 2693
rect 2693 2631 2727 2693
rect 81 97 97 2613
rect 2613 97 2629 2613
rect 2693 17 2727 79
rect -17 -17 79 17
rect 2631 -17 2727 17
<< viali >>
rect 97 97 2613 2613
<< metal1 >>
rect 85 2613 2625 2619
rect 85 97 97 2613
rect 2613 97 2625 2613
rect 85 91 2625 97
<< end >>
